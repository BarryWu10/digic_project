* SPICE NETLIST
***************************************

.SUBCKT mux21 Y A0 A1 S0 GND VDD
** N=11 EP=6 IP=0 FDC=10
* PORT Y Y 7500 52500 METAL2
* PORT A0 A0 19000 52500 METAL2
* PORT A1 A1 28000 52500 METAL2
* PORT S0 S0 39500 52500 METAL2
* PORT GND GND 26750 5000 METAL1
* PORT VDD VDD 26750 115000 METAL1
M0 8 7 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.6295e-13 $X=11500 $Y=24000 $D=1
M1 Y A0 8 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=3.564e-13 $X=17500 $Y=24000 $D=1
M2 9 A1 Y GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.346e-13 $X=25500 $Y=24000 $D=1
M3 GND S0 9 GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=3.564e-13 $X=31500 $Y=24000 $D=1
M4 7 S0 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=40000 $Y=30000 $D=1
M5 10 7 VDD VDD P L=1.8e-07 W=1.98e-06 AD=7.128e-13 AS=9.9225e-13 $X=11500 $Y=73000 $D=0
M6 Y A1 10 VDD P L=1.8e-07 W=1.98e-06 AD=1.0692e-12 AS=7.128e-13 $X=17500 $Y=73000 $D=0
M7 11 A0 Y VDD P L=1.8e-07 W=1.98e-06 AD=7.128e-13 AS=1.0692e-12 $X=25500 $Y=73000 $D=0
M8 VDD S0 11 VDD P L=1.8e-07 W=1.98e-06 AD=1.1421e-12 AS=7.128e-13 $X=31500 $Y=73000 $D=0
M9 7 S0 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.1421e-12 $X=40000 $Y=73000 $D=0
.ENDS
***************************************
.SUBCKT inv01 A Y GND VDD
** N=4 EP=4 IP=0 FDC=2
* PORT A A 10000 52500 METAL2
* PORT Y Y 19000 52500 METAL2
* PORT GND GND 12500 5000 METAL1
* PORT VDD VDD 12500 115000 METAL1
M0 Y A GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=2.9565e-13 $X=11500 $Y=26000 $D=1
M1 Y A VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.6295e-13 $X=11500 $Y=80000 $D=0
.ENDS
***************************************
.SUBCKT nor02ii A1 A0 Y VDD GND
** N=7 EP=5 IP=0 FDC=6
* PORT A1 A1 14000 52500 METAL2
* PORT A0 A0 23000 52500 METAL2
* PORT Y Y 33500 52500 METAL2
* PORT VDD VDD 20500 115000 METAL1
* PORT GND GND 20500 5000 METAL1
M0 GND A1 6 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.2275e-13 $X=11500 $Y=26000 $D=1
M1 Y A0 GND GND N L=1.8e-07 W=4.5e-07 AD=2.43e-13 AS=3.078e-13 $X=19500 $Y=26000 $D=1
M2 GND 6 Y GND N L=1.8e-07 W=4.5e-07 AD=2.9565e-13 AS=2.43e-13 $X=27500 $Y=26000 $D=1
M3 VDD A1 6 VDD P L=1.8e-07 W=9.9e-07 AD=9.1935e-13 AS=4.9005e-13 $X=11500 $Y=72000 $D=0
M4 7 A0 VDD VDD P L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=9.1935e-13 $X=20000 $Y=72000 $D=0
M5 Y 6 7 VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=5.508e-13 $X=26000 $Y=72000 $D=0
.ENDS
***************************************
.SUBCKT xnor2 A0 A1 Y GND VDD
** N=9 EP=5 IP=0 FDC=10
* PORT A0 A0 14000 52500 METAL2
* PORT A1 A1 36500 52500 METAL2
* PORT Y Y 56500 52500 METAL2
* PORT GND GND 31500 5000 METAL1
* PORT VDD VDD 31500 115000 METAL1
M0 8 A0 6 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=4.9005e-13 $X=11500 $Y=23000 $D=1
M1 GND A1 8 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=3.564e-13 $X=17500 $Y=23000 $D=1
M2 Y A1 7 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=4.9005e-13 $X=33500 $Y=23000 $D=1
M3 7 A0 Y GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.346e-13 $X=41500 $Y=23000 $D=1
M4 GND 6 7 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=5.346e-13 $X=49500 $Y=23000 $D=1
M5 6 A0 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.3025e-13 $X=18500 $Y=65500 $D=0
M6 VDD A1 6 VDD P L=1.8e-07 W=1.53e-06 AD=1.6362e-12 AS=8.262e-13 $X=26500 $Y=65500 $D=0
M7 9 A0 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.6362e-12 $X=35000 $Y=65500 $D=0
M8 Y A1 9 VDD P L=1.8e-07 W=2.88e-06 AD=1.52685e-12 AS=1.0368e-12 $X=41000 $Y=65500 $D=0
M9 VDD 6 Y VDD P L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=1.52685e-12 $X=49500 $Y=65500 $D=0
.ENDS
***************************************
.SUBCKT nand02 A1 A0 Y GND VDD
** N=6 EP=5 IP=0 FDC=4
* PORT A1 A1 8500 52500 METAL2
* PORT A0 A0 17500 52500 METAL2
* PORT Y Y 26500 52500 METAL2
* PORT GND GND 16500 5000 METAL1
* PORT VDD VDD 16500 115000 METAL1
M0 6 A1 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.6295e-13 $X=11500 $Y=19000 $D=1
M1 Y A0 6 GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=3.564e-13 $X=17500 $Y=19000 $D=1
M2 Y A1 VDD VDD P L=1.8e-07 W=1.35e-06 AD=7.29e-13 AS=6.9255e-13 $X=11500 $Y=86000 $D=0
M3 VDD A0 Y VDD P L=1.8e-07 W=1.35e-06 AD=6.9255e-13 AS=7.29e-13 $X=19500 $Y=86000 $D=0
.ENDS
***************************************
.SUBCKT nor03 Y A2 A1 A0 GND VDD
** N=8 EP=6 IP=0 FDC=6
* PORT Y Y 7500 52500 METAL2
* PORT A2 A2 16500 52500 METAL2
* PORT A1 A1 25500 52500 METAL2
* PORT A0 A0 34500 52500 METAL2
* PORT GND GND 20500 5000 METAL1
* PORT VDD VDD 20500 115000 METAL1
M0 Y A2 GND GND N L=1.8e-07 W=5.4e-07 AD=2.916e-13 AS=3.2805e-13 $X=11500 $Y=25000 $D=1
M1 GND A1 Y GND N L=1.8e-07 W=5.4e-07 AD=3.564e-13 AS=2.916e-13 $X=19500 $Y=25000 $D=1
M2 Y A0 GND GND N L=1.8e-07 W=5.4e-07 AD=2.5515e-13 AS=3.564e-13 $X=27500 $Y=25000 $D=1
M3 7 A2 Y VDD P L=1.8e-07 W=2.16e-06 AD=7.776e-13 AS=1.05705e-12 $X=15500 $Y=73000 $D=0
M4 8 A1 7 VDD P L=1.8e-07 W=2.16e-06 AD=7.776e-13 AS=7.776e-13 $X=21500 $Y=73000 $D=0
M5 VDD A0 8 VDD P L=1.8e-07 W=2.16e-06 AD=1.12995e-12 AS=7.776e-13 $X=27500 $Y=73000 $D=0
.ENDS
***************************************
.SUBCKT aoi21 A1 A0 B0 Y VDD GND
** N=8 EP=6 IP=0 FDC=6
* PORT A1 A1 8000 57500 METAL2
* PORT A0 A0 17000 57500 METAL2
* PORT B0 B0 26500 57500 METAL2
* PORT Y Y 35500 57500 METAL2
* PORT VDD VDD 20500 115000 METAL1
* PORT GND GND 20500 5000 METAL1
M0 8 A1 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.6295e-13 $X=11500 $Y=26000 $D=1
M1 Y A0 8 GND N L=1.8e-07 W=9.9e-07 AD=5.3055e-13 AS=3.564e-13 $X=17500 $Y=26000 $D=1
M2 GND B0 Y GND N L=1.8e-07 W=4.5e-07 AD=2.9565e-13 AS=5.3055e-13 $X=26000 $Y=32000 $D=1
M3 VDD A1 7 VDD P L=1.8e-07 W=1.53e-06 AD=8.91e-13 AS=7.5735e-13 $X=11500 $Y=76000 $D=0
M4 7 A0 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.91e-13 $X=19500 $Y=76000 $D=0
M5 Y B0 7 VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.262e-13 $X=27500 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=20
X0 1 2 3 7 8 xnor2 $T=0 0 0 0 $X=0 $Y=0
X1 4 5 6 7 8 xnor2 $T=64000 0 0 0 $X=64000 $Y=0
.ENDS
***************************************
.SUBCKT xor2 A0 A1 Y VDD GND
** N=10 EP=5 IP=0 FDC=12
* PORT A0 A0 12000 45000 METAL2
* PORT A1 A1 36500 45000 METAL2
* PORT Y Y 63500 45000 METAL2
* PORT VDD VDD 35500 115000 METAL1
* PORT VDD VDD 35750 115000 METAL1
* PORT GND GND 35500 5000 METAL1
* PORT GND GND 35750 5000 METAL1
M0 9 A0 6 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=4.9005e-13 $X=11500 $Y=19000 $D=1
M1 GND A1 9 GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=3.564e-13 $X=17500 $Y=19000 $D=1
M2 7 6 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.994e-13 $X=25500 $Y=19000 $D=1
M3 8 A1 7 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.346e-13 $X=33500 $Y=19000 $D=1
M4 7 A0 8 GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.346e-13 $X=41500 $Y=19000 $D=1
M5 Y 8 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=2.9565e-13 $X=57500 $Y=19000 $D=1
M6 6 A0 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.3025e-13 $X=12500 $Y=84000 $D=0
M7 VDD A1 6 VDD P L=1.8e-07 W=1.53e-06 AD=8.91e-13 AS=8.262e-13 $X=20500 $Y=84000 $D=0
M8 8 6 VDD VDD P L=1.8e-07 W=1.53e-06 AD=1.5633e-12 AS=8.91e-13 $X=28500 $Y=84000 $D=0
M9 10 A1 8 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.5633e-12 $X=37000 $Y=69000 $D=0
M10 VDD A0 10 VDD P L=1.8e-07 W=2.88e-06 AD=1.5876e-12 AS=1.0368e-12 $X=43000 $Y=69000 $D=0
M11 Y 8 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.5876e-12 $X=51500 $Y=69000 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=20
X0 1 2 3 4 8 9 mux21 $T=-1000 0 1 180 $X=-54500 $Y=0
X1 5 6 7 8 9 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7
** N=7 EP=7 IP=9 FDC=12
X0 1 2 6 7 inv01 $T=64000 0 0 0 $X=64000 $Y=0
X1 3 4 5 6 7 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT dffr D R CLK QB Q GND VDD
** N=23 EP=7 IP=0 FDC=34
* PORT D D 17000 52500 METAL2
* PORT R R 53000 52500 METAL2
* PORT CLK CLK 81500 52500 METAL2
* PORT QB QB 160000 52500 METAL2
* PORT Q Q 177500 52500 METAL2
* PORT GND GND 92500 5000 METAL1
* PORT GND GND 93750 5000 METAL1
* PORT VDD VDD 92500 115000 METAL1
* PORT VDD VDD 93750 115000 METAL1
M0 16 12 GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.3025e-13 $X=11500 $Y=21000 $D=1
M1 9 D 16 GND N L=1.8e-07 W=1.53e-06 AD=7.9785e-13 AS=5.508e-13 $X=17500 $Y=21000 $D=1
M2 17 10 9 GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=7.9785e-13 $X=26000 $Y=33000 $D=1
M3 GND 8 17 GND N L=1.8e-07 W=4.5e-07 AD=5.3055e-13 AS=1.62e-13 $X=32000 $Y=33000 $D=1
M4 10 9 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.3055e-13 $X=40500 $Y=27000 $D=1
M5 GND R 10 GND N L=1.8e-07 W=9.9e-07 AD=5.3055e-13 AS=5.346e-13 $X=48500 $Y=27000 $D=1
M6 11 10 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=5.3055e-13 $X=57000 $Y=33000 $D=1
M7 GND CLK 12 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=4.9005e-13 $X=78500 $Y=33000 $D=1
M8 8 12 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.346e-13 $X=86500 $Y=33000 $D=1
M9 13 12 14 GND N L=1.8e-07 W=4.5e-07 AD=7.9785e-13 AS=2.2275e-13 $X=108000 $Y=37500 $D=1
M10 18 11 13 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.9785e-13 $X=116500 $Y=25500 $D=1
M11 GND 8 18 GND N L=1.8e-07 W=1.53e-06 AD=8.7075e-13 AS=5.508e-13 $X=122500 $Y=25500 $D=1
M12 14 15 GND GND N L=1.8e-07 W=4.5e-07 AD=2.43e-13 AS=8.7075e-13 $X=131000 $Y=25500 $D=1
M13 GND R 14 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.43e-13 $X=139000 $Y=25500 $D=1
M14 15 13 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=3.078e-13 $X=147000 $Y=25500 $D=1
M15 GND 13 QB GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=4.9005e-13 $X=163500 $Y=19000 $D=1
M16 Q QB GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.994e-13 $X=171500 $Y=19000 $D=1
M17 19 8 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.46205e-12 $X=11500 $Y=69000 $D=0
M18 9 D 19 VDD P L=1.8e-07 W=2.88e-06 AD=1.42965e-12 AS=1.0368e-12 $X=17500 $Y=69000 $D=0
M19 20 10 9 VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=1.42965e-12 $X=26000 $Y=90500 $D=0
M20 VDD 12 20 VDD P L=1.8e-07 W=4.5e-07 AD=6.6015e-13 AS=1.62e-13 $X=32000 $Y=90500 $D=0
M21 21 9 VDD VDD P L=1.8e-07 W=1.35e-06 AD=4.86e-13 AS=6.6015e-13 $X=40500 $Y=80500 $D=0
M22 10 R 21 VDD P L=1.8e-07 W=1.35e-06 AD=6.1965e-13 AS=4.86e-13 $X=46500 $Y=80500 $D=0
M23 11 10 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=4.9005e-13 $X=62500 $Y=84500 $D=0
M24 VDD CLK 12 VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=78500 $Y=74000 $D=0
M25 8 12 VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=86500 $Y=74000 $D=0
M26 13 8 14 VDD P L=1.8e-07 W=4.5e-07 AD=1.4661e-12 AS=2.2275e-13 $X=108000 $Y=69000 $D=0
M27 22 11 13 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.4661e-12 $X=116500 $Y=69000 $D=0
M28 VDD 12 22 VDD P L=1.8e-07 W=2.88e-06 AD=1.6443e-12 AS=1.0368e-12 $X=122500 $Y=69000 $D=0
M29 23 15 VDD VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=1.6443e-12 $X=131000 $Y=69000 $D=0
M30 14 R 23 VDD P L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=1.62e-13 $X=137000 $Y=69000 $D=0
M31 15 13 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.6295e-13 $X=147000 $Y=90000 $D=0
M32 VDD 13 QB VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=163500 $Y=79000 $D=0
M33 Q QB VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=171500 $Y=79000 $D=0
.ENDS
***************************************
.SUBCKT and02 A0 A1 Y GND VDD
** N=7 EP=5 IP=0 FDC=6
* PORT A0 A0 9000 52500 METAL2
* PORT A1 A1 23000 52500 METAL2
* PORT Y Y 35000 52500 METAL2
* PORT GND GND 20750 5000 METAL1
* PORT VDD VDD 20750 115000 METAL1
M0 7 A0 6 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=4.9005e-13 $X=13500 $Y=28000 $D=1
M1 GND A1 7 GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=3.564e-13 $X=19500 $Y=28000 $D=1
M2 Y 6 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=28000 $Y=34000 $D=1
M3 6 A0 VDD VDD P L=1.8e-07 W=1.35e-06 AD=7.29e-13 AS=6.9255e-13 $X=11500 $Y=66000 $D=0
M4 VDD A1 6 VDD P L=1.8e-07 W=1.35e-06 AD=8.3025e-13 AS=7.29e-13 $X=19500 $Y=66000 $D=0
M5 Y 6 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=8.3025e-13 $X=28000 $Y=66000 $D=0
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=20
X0 1 2 3 4 8 9 mux21 $T=117500 0 1 180 $X=64000 $Y=0
X1 5 6 7 8 9 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7
** N=7 EP=7 IP=9 FDC=12
X0 1 2 6 7 inv01 $T=-1000 0 1 180 $X=-26000 $Y=0
X1 3 4 5 6 7 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT dffs_ni D S CLK Q GND VDD
** N=24 EP=6 IP=0 FDC=36
* PORT D D 17000 52500 METAL2
* PORT S S 68500 52500 METAL2
* PORT CLK CLK 93500 52500 METAL2
* PORT QB QB 172500 52500 METAL2<TRIVIAL>
* PORT Q Q 190500 52500 METAL2
* PORT GND GND 99000 5000 METAL1
* PORT VDD VDD 99000 115000 METAL1
M0 17 13 GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.3025e-13 $X=11500 $Y=21000 $D=1
M1 9 D 17 GND N L=1.8e-07 W=1.53e-06 AD=7.9785e-13 AS=5.508e-13 $X=17500 $Y=21000 $D=1
M2 18 10 9 GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=7.9785e-13 $X=26000 $Y=33000 $D=1
M3 GND 8 18 GND N L=1.8e-07 W=4.5e-07 AD=6.0345e-13 AS=1.62e-13 $X=32000 $Y=33000 $D=1
M4 19 9 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=6.0345e-13 $X=40500 $Y=27000 $D=1
M5 10 11 19 GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=3.564e-13 $X=46500 $Y=27000 $D=1
M6 GND S 11 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=4.9005e-13 $X=65500 $Y=33000 $D=1
M7 12 10 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.346e-13 $X=73500 $Y=33000 $D=1
M8 GND CLK 13 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=4.9005e-13 $X=90500 $Y=33000 $D=1
M9 8 13 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.346e-13 $X=98500 $Y=33000 $D=1
M10 14 13 15 GND N L=1.8e-07 W=4.5e-07 AD=7.9785e-13 AS=2.2275e-13 $X=120000 $Y=36000 $D=1
M11 20 12 14 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.9785e-13 $X=128500 $Y=24000 $D=1
M12 GND 8 20 GND N L=1.8e-07 W=1.53e-06 AD=8.7075e-13 AS=5.508e-13 $X=134500 $Y=24000 $D=1
M13 21 16 GND GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=8.7075e-13 $X=143000 $Y=36000 $D=1
M14 15 11 21 GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=1.62e-13 $X=149000 $Y=36000 $D=1
M15 16 14 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=2.9565e-13 $X=159500 $Y=19000 $D=1
M16 GND 14 QB GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=4.9005e-13 $X=176500 $Y=19000 $D=1
M17 Q QB GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.994e-13 $X=184500 $Y=19000 $D=1
M18 22 8 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.46205e-12 $X=11500 $Y=69000 $D=0
M19 9 D 22 VDD P L=1.8e-07 W=2.88e-06 AD=1.42965e-12 AS=1.0368e-12 $X=17500 $Y=69000 $D=0
M20 23 10 9 VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=1.42965e-12 $X=26000 $Y=90500 $D=0
M21 VDD 13 23 VDD P L=1.8e-07 W=4.5e-07 AD=6.6015e-13 AS=1.62e-13 $X=32000 $Y=90500 $D=0
M22 10 9 VDD VDD P L=1.8e-07 W=1.35e-06 AD=7.29e-13 AS=6.6015e-13 $X=40500 $Y=80500 $D=0
M23 VDD 11 10 VDD P L=1.8e-07 W=1.35e-06 AD=6.1965e-13 AS=7.29e-13 $X=48500 $Y=80500 $D=0
M24 VDD S 11 VDD P L=1.8e-07 W=1.98e-06 AD=1.0692e-12 AS=9.1935e-13 $X=65500 $Y=74000 $D=0
M25 12 10 VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.0692e-12 $X=73500 $Y=74000 $D=0
M26 VDD CLK 13 VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=90500 $Y=74000 $D=0
M27 8 13 VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=98500 $Y=74000 $D=0
M28 14 8 15 VDD P L=1.8e-07 W=4.5e-07 AD=1.4661e-12 AS=2.2275e-13 $X=120000 $Y=69000 $D=0
M29 24 12 14 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.4661e-12 $X=128500 $Y=69000 $D=0
M30 VDD 13 24 VDD P L=1.8e-07 W=2.88e-06 AD=1.60785e-12 AS=1.0368e-12 $X=134500 $Y=69000 $D=0
M31 15 16 VDD VDD P L=1.8e-07 W=4.5e-07 AD=2.43e-13 AS=1.60785e-12 $X=143000 $Y=79000 $D=0
M32 VDD 11 15 VDD P L=1.8e-07 W=4.5e-07 AD=6.0345e-13 AS=2.43e-13 $X=151000 $Y=79000 $D=0
M33 16 14 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=6.0345e-13 $X=159500 $Y=73000 $D=0
M34 VDD 14 QB VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=176500 $Y=79000 $D=0
M35 Q QB VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=184500 $Y=79000 $D=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=20
X0 1 2 3 4 8 9 mux21 $T=64000 0 0 0 $X=64000 $Y=0
X1 5 6 7 8 9 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT and03 A0 A1 A2 Y GND VDD
** N=9 EP=6 IP=0 FDC=8
* PORT A0 A0 11500 52500 METAL2
* PORT A1 A1 20500 52500 METAL2
* PORT A2 A2 29500 52500 METAL2
* PORT Y Y 42500 52500 METAL2
* PORT GND GND 24750 5000 METAL1
* PORT VDD VDD 24750 115000 METAL1
M0 8 A0 7 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.5735e-13 $X=13500 $Y=26000 $D=1
M1 9 A1 8 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=5.508e-13 $X=19500 $Y=26000 $D=1
M2 GND A2 9 GND N L=1.8e-07 W=1.53e-06 AD=8.7075e-13 AS=5.508e-13 $X=25500 $Y=26000 $D=1
M3 Y 7 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=8.7075e-13 $X=34000 $Y=38000 $D=1
M4 VDD A0 7 VDD P L=1.8e-07 W=1.8e-06 AD=1.0368e-12 AS=8.5455e-13 $X=11500 $Y=72000 $D=0
M5 7 A1 VDD VDD P L=1.8e-07 W=1.8e-06 AD=9.72e-13 AS=1.0368e-12 $X=19500 $Y=72000 $D=0
M6 VDD A2 7 VDD P L=1.8e-07 W=1.8e-06 AD=1.053e-12 AS=9.72e-13 $X=27500 $Y=72000 $D=0
M7 Y 7 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.053e-12 $X=36000 $Y=72000 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=20
X0 1 2 3 7 8 xnor2 $T=0 0 0 0 $X=0 $Y=0
X1 4 5 6 7 8 xnor2 $T=127000 0 1 180 $X=64000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=30
X0 1 2 3 4 11 12 mux21 $T=128000 0 0 0 $X=128000 $Y=0
X1 5 6 7 10 9 8 11 12 ICV_7 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=20
X0 1 2 3 7 8 xnor2 $T=-64000 0 0 0 $X=-64000 $Y=0
X1 4 5 6 7 8 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=16
X0 1 2 3 8 7 nor02ii $T=-1000 0 1 180 $X=-42000 $Y=0
X1 4 5 6 7 8 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT and04 A0 A1 A2 A3 Y GND VDD
** N=11 EP=7 IP=0 FDC=10
* PORT A0 A0 12000 52500 METAL2
* PORT A1 A1 21000 52500 METAL2
* PORT A2 A2 30000 52500 METAL2
* PORT A3 A3 39000 52500 METAL2
* PORT Y Y 51000 52500 METAL2
* PORT GND GND 28750 5000 METAL1
* PORT VDD VDD 28750 115000 METAL1
M0 9 A0 8 GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=1.02465e-12 $X=15500 $Y=20000 $D=1
M1 10 A1 9 GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=7.452e-13 $X=21500 $Y=20000 $D=1
M2 11 A2 10 GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=7.452e-13 $X=27500 $Y=20000 $D=1
M3 GND A3 11 GND N L=1.8e-07 W=2.07e-06 AD=1.13805e-12 AS=7.452e-13 $X=33500 $Y=20000 $D=1
M4 Y 8 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=1.13805e-12 $X=42000 $Y=38000 $D=1
M5 8 A0 VDD VDD P L=1.8e-07 W=2.25e-06 AD=1.215e-12 AS=1.16235e-12 $X=11500 $Y=69500 $D=0
M6 VDD A1 8 VDD P L=1.8e-07 W=2.25e-06 AD=1.2798e-12 AS=1.215e-12 $X=19500 $Y=69500 $D=0
M7 8 A2 VDD VDD P L=1.8e-07 W=2.25e-06 AD=1.215e-12 AS=1.2798e-12 $X=27500 $Y=69500 $D=0
M8 VDD A3 8 VDD P L=1.8e-07 W=2.25e-06 AD=1.27575e-12 AS=1.215e-12 $X=35500 $Y=69500 $D=0
M9 Y 8 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.27575e-12 $X=44000 $Y=69500 $D=0
.ENDS
***************************************
.SUBCKT aoi22 Y B1 B0 A0 A1 VDD GND
** N=10 EP=7 IP=0 FDC=8
* PORT Y Y 6500 52500 METAL2
* PORT B1 B1 15500 52500 METAL2
* PORT B0 B0 24500 52500 METAL2
* PORT A0 A0 33500 52500 METAL2
* PORT A1 A1 42500 52500 METAL2
* PORT VDD VDD 24500 115000 METAL1
* PORT GND GND 24500 5000 METAL1
M0 9 B1 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.6295e-13 $X=13500 $Y=26000 $D=1
M1 Y B0 9 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=3.564e-13 $X=19500 $Y=26000 $D=1
M2 10 A0 Y GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.346e-13 $X=27500 $Y=26000 $D=1
M3 GND A1 10 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=3.564e-13 $X=33500 $Y=26000 $D=1
M4 Y B1 8 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=7.5735e-13 $X=11500 $Y=72000 $D=0
M5 8 B0 Y VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=19500 $Y=72000 $D=0
M6 VDD A0 8 VDD P L=1.8e-07 W=1.53e-06 AD=8.91e-13 AS=8.262e-13 $X=27500 $Y=72000 $D=0
M7 8 A1 VDD VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.91e-13 $X=35500 $Y=72000 $D=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=30
X0 1 2 3 4 11 12 mux21 $T=-65000 0 1 180 $X=-118500 $Y=0
X1 5 6 7 8 9 10 11 12 ICV_9 $T=0 0 0 0 $X=-64000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=20
X0 1 2 3 4 8 9 mux21 $T=-54500 0 0 0 $X=-54500 $Y=0
X1 5 6 7 8 9 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT nand04 A0 Y A1 A2 A3 GND VDD
** N=10 EP=7 IP=0 FDC=8
* PORT A0 A0 6500 60000 METAL2
* PORT Y Y 15500 60000 METAL2
* PORT A1 A1 24500 60000 METAL2
* PORT A2 A2 33500 60000 METAL2
* PORT A3 A3 42500 60000 METAL2
* PORT GND GND 24500 5000 METAL1
* PORT VDD VDD 24500 115000 METAL1
M0 8 A0 Y GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=1.02465e-12 $X=14500 $Y=21000 $D=1
M1 9 A1 8 GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=7.452e-13 $X=20500 $Y=21000 $D=1
M2 10 A2 9 GND N L=1.8e-07 W=2.07e-06 AD=7.452e-13 AS=7.452e-13 $X=26500 $Y=21000 $D=1
M3 GND A3 10 GND N L=1.8e-07 W=2.07e-06 AD=1.09755e-12 AS=7.452e-13 $X=32500 $Y=21000 $D=1
M4 Y A0 VDD VDD P L=1.8e-07 W=2.16e-06 AD=1.1664e-12 AS=1.12995e-12 $X=11500 $Y=75000 $D=0
M5 VDD A1 Y VDD P L=1.8e-07 W=2.16e-06 AD=1.2312e-12 AS=1.1664e-12 $X=19500 $Y=75000 $D=0
M6 Y A2 VDD VDD P L=1.8e-07 W=2.16e-06 AD=1.1664e-12 AS=1.2312e-12 $X=27500 $Y=75000 $D=0
M7 VDD A3 Y VDD P L=1.8e-07 W=2.16e-06 AD=1.12995e-12 AS=1.1664e-12 $X=35500 $Y=75000 $D=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=30
X0 1 2 3 4 11 12 mux21 $T=181500 0 1 180 $X=128000 $Y=0
X1 5 6 7 10 9 8 11 12 ICV_7 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT mux21_ni S0 A1 A0 Y GND VDD
** N=12 EP=6 IP=0 FDC=12
* PORT S0 S0 14500 52500 METAL2
* PORT A1 A1 24500 52500 METAL2
* PORT A0 A0 33500 52500 METAL2
* PORT Y Y 55500 52500 METAL2
* PORT GND GND 31000 5000 METAL1
* PORT VDD VDD 31000 115000 METAL1
M0 GND S0 7 GND N L=1.8e-07 W=4.5e-07 AD=6.0345e-13 AS=2.2275e-13 $X=11500 $Y=27500 $D=1
M1 9 S0 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=6.0345e-13 $X=20000 $Y=21500 $D=1
M2 8 A1 9 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=3.564e-13 $X=26000 $Y=21500 $D=1
M3 10 A0 8 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.346e-13 $X=34000 $Y=21500 $D=1
M4 GND 7 10 GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=3.564e-13 $X=40000 $Y=21500 $D=1
M5 Y 8 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=48500 $Y=27500 $D=1
M6 VDD S0 7 VDD P L=1.8e-07 W=9.9e-07 AD=1.1421e-12 AS=4.9005e-13 $X=11500 $Y=78000 $D=0
M7 11 S0 VDD VDD P L=1.8e-07 W=1.98e-06 AD=7.128e-13 AS=1.1421e-12 $X=20000 $Y=78000 $D=0
M8 8 A0 11 VDD P L=1.8e-07 W=1.98e-06 AD=1.0692e-12 AS=7.128e-13 $X=26000 $Y=78000 $D=0
M9 12 A1 8 VDD P L=1.8e-07 W=1.98e-06 AD=7.128e-13 AS=1.0692e-12 $X=34000 $Y=78000 $D=0
M10 VDD 7 12 VDD P L=1.8e-07 W=1.98e-06 AD=1.1421e-12 AS=7.128e-13 $X=40000 $Y=78000 $D=0
M11 Y 8 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.1421e-12 $X=48500 $Y=78000 $D=0
.ENDS
***************************************
.SUBCKT latchr CLK D R QB GND VDD
** N=14 EP=6 IP=0 FDC=16
* PORT CLK CLK 14500 52500 METAL2
* PORT D D 27500 52500 METAL2
* PORT R R 57500 52500 METAL2
* PORT QB QB 76500 52500 METAL2
* PORT GND GND 42500 5000 METAL1
* PORT VDD VDD 42500 115000 METAL1
M0 GND CLK 7 GND N L=1.8e-07 W=4.5e-07 AD=8.7075e-13 AS=2.2275e-13 $X=11500 $Y=33000 $D=1
M1 10 CLK GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.7075e-13 $X=20000 $Y=21000 $D=1
M2 8 D 10 GND N L=1.8e-07 W=1.53e-06 AD=7.9785e-13 AS=5.508e-13 $X=26000 $Y=21000 $D=1
M3 11 7 8 GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=7.9785e-13 $X=34500 $Y=25000 $D=1
M4 GND 9 11 GND N L=1.8e-07 W=4.5e-07 AD=6.0345e-13 AS=1.62e-13 $X=40500 $Y=25000 $D=1
M5 9 8 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=6.0345e-13 $X=49000 $Y=19000 $D=1
M6 GND R 9 GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=5.346e-13 $X=57000 $Y=19000 $D=1
M7 QB 9 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=65500 $Y=25000 $D=1
M8 VDD CLK 7 VDD P L=1.8e-07 W=9.9e-07 AD=1.5876e-12 AS=4.9005e-13 $X=11500 $Y=69000 $D=0
M9 12 7 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.5876e-12 $X=20000 $Y=69000 $D=0
M10 8 D 12 VDD P L=1.8e-07 W=2.88e-06 AD=1.42965e-12 AS=1.0368e-12 $X=26000 $Y=69000 $D=0
M11 13 CLK 8 VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=1.42965e-12 $X=34500 $Y=83000 $D=0
M12 VDD 9 13 VDD P L=1.8e-07 W=4.5e-07 AD=9.153e-13 AS=1.62e-13 $X=40500 $Y=83000 $D=0
M13 14 8 VDD VDD P L=1.8e-07 W=1.62e-06 AD=5.832e-13 AS=9.153e-13 $X=49000 $Y=83000 $D=0
M14 9 R 14 VDD P L=1.8e-07 W=1.62e-06 AD=7.8975e-13 AS=5.832e-13 $X=55000 $Y=83000 $D=0
M15 QB 9 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.6295e-13 $X=71500 $Y=90000 $D=0
.ENDS
***************************************
.SUBCKT oai22 A0 A1 Y B1 B0 GND VDD
** N=10 EP=7 IP=0 FDC=8
* PORT A0 A0 6500 52500 METAL2
* PORT A1 A1 15500 52500 METAL2
* PORT Y Y 24500 52500 METAL2
* PORT B1 B1 33500 52500 METAL2
* PORT B0 B0 42500 52500 METAL2
* PORT GND GND 24500 5000 METAL1
* PORT VDD VDD 24500 115000 METAL1
M0 Y A0 8 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=4.9005e-13 $X=11500 $Y=22500 $D=1
M1 8 A1 Y GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.346e-13 $X=19500 $Y=22500 $D=1
M2 GND B1 8 GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=5.346e-13 $X=27500 $Y=22500 $D=1
M3 8 B0 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.994e-13 $X=35500 $Y=22500 $D=1
M4 9 A0 VDD VDD P L=1.8e-07 W=2.61e-06 AD=9.396e-13 AS=1.36485e-12 $X=13500 $Y=66000 $D=0
M5 Y A1 9 VDD P L=1.8e-07 W=2.61e-06 AD=1.4094e-12 AS=9.396e-13 $X=19500 $Y=66000 $D=0
M6 10 B1 Y VDD P L=1.8e-07 W=2.61e-06 AD=9.396e-13 AS=1.4094e-12 $X=27500 $Y=66000 $D=0
M7 VDD B0 10 VDD P L=1.8e-07 W=2.61e-06 AD=1.36485e-12 AS=9.396e-13 $X=33500 $Y=66000 $D=0
.ENDS
***************************************
.SUBCKT oai21 B0 A1 Y A0 GND VDD
** N=8 EP=6 IP=0 FDC=6
* PORT B0 B0 6500 52500 METAL2
* PORT A1 A1 15500 52500 METAL2
* PORT Y Y 24500 52500 METAL2
* PORT A0 A0 33500 52500 METAL2
* PORT GND GND 20500 5000 METAL1
* PORT VDD VDD 20500 115000 METAL1
M0 7 B0 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.6295e-13 $X=11500 $Y=25000 $D=1
M1 Y A1 7 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.346e-13 $X=19500 $Y=25000 $D=1
M2 7 A0 Y GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.346e-13 $X=27500 $Y=25000 $D=1
M3 Y B0 VDD VDD P L=1.8e-07 W=1.35e-06 AD=1.41345e-12 AS=6.9255e-13 $X=13000 $Y=68000 $D=0
M4 8 A1 Y VDD P L=1.8e-07 W=2.61e-06 AD=9.396e-13 AS=1.41345e-12 $X=21500 $Y=68000 $D=0
M5 VDD A0 8 VDD P L=1.8e-07 W=2.61e-06 AD=1.36485e-12 AS=9.396e-13 $X=27500 $Y=68000 $D=0
.ENDS
***************************************
.SUBCKT nor02 A1 Y A0 VDD GND
** N=6 EP=5 IP=0 FDC=4
* PORT A1 A1 7500 57500 METAL2
* PORT Y Y 16500 57500 METAL2
* PORT A0 A0 25500 57500 METAL2
* PORT VDD VDD 16500 115000 METAL1
* PORT GND GND 16500 5000 METAL1
M0 Y A1 GND GND N L=1.8e-07 W=4.5e-07 AD=2.43e-13 AS=2.9565e-13 $X=11500 $Y=26000 $D=1
M1 GND A0 Y GND N L=1.8e-07 W=4.5e-07 AD=2.9565e-13 AS=2.43e-13 $X=19500 $Y=26000 $D=1
M2 6 A1 Y VDD P L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.5735e-13 $X=11500 $Y=76000 $D=0
M3 VDD A0 6 VDD P L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=5.508e-13 $X=17500 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT or02 A1 A0 Y VDD GND
** N=7 EP=5 IP=0 FDC=6
* PORT A1 A1 12500 52500 METAL2
* PORT A0 A0 21500 52500 METAL2
* PORT Y Y 33500 52500 METAL2
* PORT VDD VDD 20500 115000 METAL1
* PORT GND GND 20500 5000 METAL1
M0 6 A1 GND GND N L=1.8e-07 W=4.5e-07 AD=2.43e-13 AS=2.9565e-13 $X=11500 $Y=19000 $D=1
M1 GND A0 6 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.43e-13 $X=19500 $Y=19000 $D=1
M2 Y 6 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=3.078e-13 $X=27500 $Y=19000 $D=1
M3 7 A1 6 VDD P L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.5735e-13 $X=13000 $Y=84000 $D=0
M4 VDD A0 7 VDD P L=1.8e-07 W=1.53e-06 AD=9.1935e-13 AS=5.508e-13 $X=19000 $Y=84000 $D=0
M5 Y 6 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=9.1935e-13 $X=27500 $Y=84000 $D=0
.ENDS
***************************************
.SUBCKT aoi32 A2 A1 A0 Y B0 B1 VDD GND
** N=12 EP=8 IP=0 FDC=10
* PORT A2 A2 5500 52500 METAL2
* PORT A1 A1 14500 52500 METAL2
* PORT A0 A0 23500 52500 METAL2
* PORT Y Y 32500 52500 METAL2
* PORT B0 B0 41500 52500 METAL2
* PORT B1 B1 50500 52500 METAL2
* PORT VDD VDD 28500 115000 METAL1
* PORT GND GND 28500 5000 METAL1
M0 10 A2 GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.3025e-13 $X=11500 $Y=19500 $D=1
M1 11 A1 10 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=5.508e-13 $X=17500 $Y=19500 $D=1
M2 Y A0 11 GND N L=1.8e-07 W=1.53e-06 AD=8.4645e-13 AS=5.508e-13 $X=23500 $Y=19500 $D=1
M3 12 B0 Y GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=8.4645e-13 $X=32000 $Y=25500 $D=1
M4 GND B1 12 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=3.564e-13 $X=38000 $Y=25500 $D=1
M5 9 A2 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.3025e-13 $X=11500 $Y=81000 $D=0
M6 VDD A1 9 VDD P L=1.8e-07 W=1.53e-06 AD=8.91e-13 AS=8.262e-13 $X=19500 $Y=81000 $D=0
M7 9 A0 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.91e-13 $X=27500 $Y=81000 $D=0
M8 Y B0 9 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=35500 $Y=81000 $D=0
M9 9 B1 Y VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.262e-13 $X=43500 $Y=81000 $D=0
.ENDS
***************************************
.SUBCKT nand03 A0 Y A1 A2 VDD GND
** N=8 EP=6 IP=0 FDC=6
* PORT A0 A0 7500 55000 METAL2
* PORT Y Y 16500 55000 METAL2
* PORT A1 A1 25500 55000 METAL2
* PORT A2 A2 34500 55000 METAL2
* PORT VDD VDD 20500 115000 METAL1
* PORT GND GND 20500 5000 METAL1
M0 7 A0 Y GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.5735e-13 $X=13500 $Y=24500 $D=1
M1 8 A1 7 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=5.508e-13 $X=19500 $Y=24500 $D=1
M2 GND A2 8 GND N L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=5.508e-13 $X=25500 $Y=24500 $D=1
M3 Y A0 VDD VDD P L=1.8e-07 W=1.62e-06 AD=8.748e-13 AS=8.6265e-13 $X=11500 $Y=74000 $D=0
M4 VDD A1 Y VDD P L=1.8e-07 W=1.62e-06 AD=9.396e-13 AS=8.748e-13 $X=19500 $Y=74000 $D=0
M5 Y A2 VDD VDD P L=1.8e-07 W=1.62e-06 AD=7.8975e-13 AS=9.396e-13 $X=27500 $Y=74000 $D=0
.ENDS
***************************************
.SUBCKT aoi221 C0 B0 B1 Y A1 A0 GND VDD
** N=12 EP=8 IP=0 FDC=10
* PORT C0 C0 9500 52500 METAL2
* PORT B0 B0 18500 52500 METAL2
* PORT B1 B1 27500 52500 METAL2
* PORT Y Y 36500 52500 METAL2
* PORT A1 A1 45500 52500 METAL2
* PORT A0 A0 54500 52500 METAL2
* PORT GND GND 32500 5000 METAL1
* PORT VDD VDD 32500 115000 METAL1
M0 Y C0 GND GND N L=1.8e-07 W=4.5e-07 AD=5.3055e-13 AS=2.9565e-13 $X=11500 $Y=32000 $D=1
M1 11 B0 Y GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.3055e-13 $X=20000 $Y=26000 $D=1
M2 GND B1 11 GND N L=1.8e-07 W=9.9e-07 AD=7.4115e-13 AS=3.564e-13 $X=26000 $Y=26000 $D=1
M3 12 A1 GND GND N L=1.8e-07 W=1.17e-06 AD=4.212e-13 AS=7.4115e-13 $X=34500 $Y=24000 $D=1
M4 Y A0 12 GND N L=1.8e-07 W=1.17e-06 AD=5.5485e-13 AS=4.212e-13 $X=40500 $Y=24000 $D=1
M5 9 C0 Y VDD P L=1.8e-07 W=2.07e-06 AD=1.1178e-12 AS=1.02465e-12 $X=11500 $Y=73000 $D=0
M6 10 B0 9 VDD P L=1.8e-07 W=2.07e-06 AD=1.1178e-12 AS=1.1178e-12 $X=19500 $Y=73000 $D=0
M7 9 B1 10 VDD P L=1.8e-07 W=2.07e-06 AD=1.02465e-12 AS=1.1178e-12 $X=27500 $Y=73000 $D=0
M8 VDD A1 10 VDD P L=1.8e-07 W=2.07e-06 AD=1.1826e-12 AS=1.02465e-12 $X=43500 $Y=73000 $D=0
M9 10 A0 VDD VDD P L=1.8e-07 W=2.07e-06 AD=1.02465e-12 AS=1.1826e-12 $X=51500 $Y=73000 $D=0
.ENDS
***************************************
.SUBCKT ao22 A1 A0 B0 B1 Y GND VDD
** N=11 EP=7 IP=0 FDC=10
* PORT A1 A1 6000 52500 METAL2
* PORT A0 A0 15000 52500 METAL2
* PORT B0 B0 24000 52500 METAL2
* PORT B1 B1 34000 52500 METAL2
* PORT Y Y 51000 52500 METAL2
* PORT GND GND 28750 5000 METAL1
* PORT VDD VDD 28750 115000 METAL1
M0 10 A1 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.6295e-13 $X=13500 $Y=26000 $D=1
M1 9 A0 10 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=3.564e-13 $X=19500 $Y=26000 $D=1
M2 11 B0 9 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.346e-13 $X=27500 $Y=26000 $D=1
M3 GND B1 11 GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=3.564e-13 $X=33500 $Y=26000 $D=1
M4 Y 9 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=42000 $Y=32000 $D=1
M5 8 A1 VDD VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.3025e-13 $X=11500 $Y=72000 $D=0
M6 9 B0 8 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=19500 $Y=72000 $D=0
M7 8 B1 9 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=27500 $Y=72000 $D=0
M8 VDD A0 8 VDD P L=1.8e-07 W=1.53e-06 AD=9.1935e-13 AS=8.262e-13 $X=35500 $Y=72000 $D=0
M9 Y 9 VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=9.1935e-13 $X=44000 $Y=72000 $D=0
.ENDS
***************************************
.SUBCKT buf02 Y A GND VDD
** N=5 EP=4 IP=0 FDC=4
* PORT Y Y 7500 52500 METAL2
* PORT A A 19500 52500 METAL2
* PORT GND GND 16750 5000 METAL1
* PORT VDD VDD 16750 115000 METAL1
M0 GND 5 Y GND N L=1.8e-07 W=9.9e-07 AD=6.0345e-13 AS=4.9005e-13 $X=11500 $Y=25000 $D=1
M1 5 A GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=6.0345e-13 $X=20000 $Y=31000 $D=1
M2 VDD 5 Y VDD P L=1.8e-07 W=1.98e-06 AD=1.1421e-12 AS=9.1935e-13 $X=11500 $Y=71000 $D=0
M3 5 A VDD VDD P L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=1.1421e-12 $X=20000 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT sobel_layout o_mode[1] i_reset i_pixel_bot[16] i_pixel_bot[0] i_pixel_top[15] i_pixel_mid[17] i_pixel_bot[7] i_pixel_mid[7] i_pixel_bot[2] i_pixel_top[1] i_clock i_pixel_mid[16] i_pixel_top[17] i_pixel_bot[9] i_valid i_pixel_top[16] i_pixel_bot[18] i_pixel_top[19] i_pixel_top[0] i_pixel_top[11]
+ i_pixel_mid[22] i_pixel_top[9] i_pixel_mid[0] i_pixel_bot[3] i_pixel_mid[3] i_pixel_mid[2] i_pixel_mid[18] i_pixel_top[3] i_pixel_bot[14] i_pixel_bot[11] i_pixel_bot[6] o_mode[0] i_pixel_bot[4] i_pixel_top[21] i_pixel_bot[19] i_pixel_mid[4] i_pixel_bot[13] i_pixel_bot[12] i_pixel_top[4] i_pixel_top[5]
+ i_pixel_mid[20] i_pixel_bot[20] i_pixel_bot[21] i_pixel_mid[5] i_pixel_bot[15] i_pixel_top[7] i_pixel_top[20] i_pixel_mid[23] i_pixel_top[12] i_pixel_top[13] o_dir[0] i_pixel_bot[1] i_pixel_bot[8] i_pixel_top[8] i_pixel_top[18] i_pixel_mid[1] i_pixel_bot[17] i_pixel_top[2] o_dir[2] o_valid
+ o_dir[1] o_edge i_pixel_mid[21] i_pixel_mid[19] i_pixel_top[22] i_pixel_bot[5] i_pixel_mid[6] i_pixel_bot[22] i_pixel_bot[10] i_pixel_top[6] i_pixel_top[23] i_pixel_top[14] i_pixel_bot[23] i_pixel_top[10] VDD GND
** N=1363 EP=76 IP=5964 FDC=11184
* PORT o_mode[1] o_mode[1] 5500 1121000 METAL5
* PORT i_reset i_reset 5500 1706000 METAL5
* PORT i_pixel_bot[16] i_pixel_bot[16] 5500 1686000 METAL5
* PORT i_pixel_bot[0] i_pixel_bot[0] 5500 1696000 METAL5
* PORT i_pixel_top[15] i_pixel_top[15] 5500 1616000 METAL5
* PORT i_pixel_mid[17] i_pixel_mid[17] 5500 1676000 METAL5
* PORT i_pixel_bot[7] i_pixel_bot[7] 5500 1566000 METAL5
* PORT i_pixel_mid[7] i_pixel_mid[7] 5500 1576000 METAL5
* PORT i_pixel_bot[2] i_pixel_bot[2] 5500 1646000 METAL5
* PORT i_pixel_top[1] i_pixel_top[1] 5500 1656000 METAL5
* PORT i_clock i_clock 2122000 2500 METAL4
* PORT i_pixel_mid[16] i_pixel_mid[16] 3842500 1682000 METAL5
* PORT i_pixel_top[17] i_pixel_top[17] 3842500 1692000 METAL5
* PORT i_pixel_bot[9] i_pixel_bot[9] 2100000 3053000 METAL4
* PORT i_valid i_valid 3842500 1712000 METAL5
* PORT i_pixel_top[16] i_pixel_top[16] 2100000 2500 METAL4
* PORT i_pixel_bot[18] i_pixel_bot[18] 5500 1586000 METAL5
* PORT i_pixel_top[19] i_pixel_top[19] 5500 1636000 METAL5
* PORT i_pixel_top[0] i_pixel_top[0] 3842500 1702000 METAL5
* PORT i_pixel_top[11] i_pixel_top[11] 5500 1626000 METAL5
* PORT i_pixel_mid[22] i_pixel_mid[22] 5500 1546000 METAL5
* PORT i_pixel_top[9] i_pixel_top[9] 5500 1666000 METAL5
* PORT i_pixel_mid[0] i_pixel_mid[0] 2122000 3053000 METAL4
* PORT i_pixel_bot[3] i_pixel_bot[3] 3842500 1575000 METAL5
* PORT i_pixel_mid[3] i_pixel_mid[3] 1946000 2500 METAL4
* PORT i_pixel_mid[2] i_pixel_mid[2] 3842500 1635000 METAL5
* PORT i_pixel_mid[18] i_pixel_mid[18] 2023000 3053000 METAL4
* PORT i_pixel_top[3] i_pixel_top[3] 1968000 2500 METAL4
* PORT i_pixel_bot[14] i_pixel_bot[14] 1957000 2500 METAL4
* PORT i_pixel_bot[11] i_pixel_bot[11] 3842500 1615000 METAL5
* PORT i_pixel_bot[6] i_pixel_bot[6] 2034000 3053000 METAL4
* PORT o_mode[0] o_mode[0] 1946000 3053000 METAL4
* PORT i_pixel_bot[4] i_pixel_bot[4] 2034000 2500 METAL4
* PORT i_pixel_top[21] i_pixel_top[21] 2045000 2500 METAL4
* PORT i_pixel_bot[19] i_pixel_bot[19] 2067000 2500 METAL4
* PORT i_pixel_mid[4] i_pixel_mid[4] 1990000 2500 METAL4
* PORT i_pixel_bot[13] i_pixel_bot[13] 2012000 2500 METAL4
* PORT i_pixel_bot[12] i_pixel_bot[12] 3842500 1565000 METAL5
* PORT i_pixel_top[4] i_pixel_top[4] 5500 1606000 METAL5
* PORT i_pixel_top[5] i_pixel_top[5] 5500 1556000 METAL5
* PORT i_pixel_mid[20] i_pixel_mid[20] 3842500 1555000 METAL5
* PORT i_pixel_bot[20] i_pixel_bot[20] 3842500 1605000 METAL5
* PORT i_pixel_bot[21] i_pixel_bot[21] 3842500 1655000 METAL5
* PORT i_pixel_mid[5] i_pixel_mid[5] 3842500 1545000 METAL5
* PORT i_pixel_bot[15] i_pixel_bot[15] 5500 1596000 METAL5
* PORT i_pixel_top[7] i_pixel_top[7] 3842500 1595000 METAL5
* PORT i_pixel_top[20] i_pixel_top[20] 3842500 1585000 METAL5
* PORT i_pixel_mid[23] i_pixel_mid[23] 3842500 1645000 METAL5
* PORT i_pixel_top[12] i_pixel_top[12] 3842500 1665000 METAL5
* PORT i_pixel_top[13] i_pixel_top[13] 3842500 1625000 METAL5
* PORT o_dir[0] o_dir[0] 3842500 1450000 METAL5
* PORT i_pixel_bot[1] i_pixel_bot[1] 2056000 2500 METAL4
* PORT i_pixel_bot[8] i_pixel_bot[8] 2111000 3053000 METAL4
* PORT i_pixel_top[8] i_pixel_top[8] 2111000 2500 METAL4
* PORT i_pixel_top[18] i_pixel_top[18] 2056000 3053000 METAL4
* PORT i_pixel_mid[1] i_pixel_mid[1] 2089000 3053000 METAL4
* PORT i_pixel_bot[17] i_pixel_bot[17] 2089000 2500 METAL4
* PORT i_pixel_top[2] i_pixel_top[2] 2023000 2500 METAL4
* PORT o_dir[2] o_dir[2] 1924000 2500 METAL4
* PORT o_valid o_valid 1924000 3053000 METAL4
* PORT o_dir[1] o_dir[1] 1935000 3053000 METAL4
* PORT o_edge o_edge 1935000 2500 METAL4
* PORT i_pixel_mid[21] i_pixel_mid[21] 1957000 3053000 METAL4
* PORT i_pixel_mid[19] i_pixel_mid[19] 1968000 3053000 METAL4
* PORT i_pixel_top[22] i_pixel_top[22] 1979000 2500 METAL4
* PORT i_pixel_bot[5] i_pixel_bot[5] 1979000 3053000 METAL4
* PORT i_pixel_mid[6] i_pixel_mid[6] 1990000 3053000 METAL4
* PORT i_pixel_bot[22] i_pixel_bot[22] 2001000 2500 METAL4
* PORT i_pixel_bot[10] i_pixel_bot[10] 2001000 3053000 METAL4
* PORT i_pixel_top[6] i_pixel_top[6] 2012000 3053000 METAL4
* PORT i_pixel_top[23] i_pixel_top[23] 2045000 3053000 METAL4
* PORT i_pixel_top[14] i_pixel_top[14] 2078000 3053000 METAL4
* PORT i_pixel_bot[23] i_pixel_bot[23] 2067000 3053000 METAL4
* PORT i_pixel_top[10] i_pixel_top[10] 2078000 2500 METAL4
* PORT VDD VDD 3842500 1416500 METAL1
* PORT GND GND 5500 1087500 METAL1
M0 404 1299 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.6295e-13 $X=163500 $Y=172500 $D=1
M1 GND 406 404 GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=5.346e-13 $X=171500 $Y=172500 $D=1
M2 404 417 GND GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=5.994e-13 $X=179500 $Y=172500 $D=1
M3 GND 422 404 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=5.346e-13 $X=187500 $Y=172500 $D=1
M4 1329 535 539 GND N L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=7.5735e-13 $X=723500 $Y=935000 $D=1
M5 539 575 1329 GND N L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=731500 $Y=935000 $D=1
M6 1329 31 539 GND N L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.262e-13 $X=739500 $Y=935000 $D=1
M7 1329 199 1330 GND N L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=7.5735e-13 $X=755500 $Y=935000 $D=1
M8 1330 194 1329 GND N L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=763500 $Y=935000 $D=1
M9 GND 584 1330 GND N L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=8.262e-13 $X=771500 $Y=935000 $D=1
M10 GND 1331 659 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.2275e-13 $X=963500 $Y=954000 $D=1
M11 1331 224 GND GND N L=1.8e-07 W=4.5e-07 AD=5.3055e-13 AS=3.078e-13 $X=971500 $Y=954000 $D=1
M12 1342 649 1331 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.3055e-13 $X=980000 $Y=948000 $D=1
M13 GND 205 1342 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=3.564e-13 $X=986000 $Y=948000 $D=1
M14 1343 265 741 GND N L=1.8e-07 W=1.17e-06 AD=4.212e-13 AS=5.5485e-13 $X=1379500 $Y=940500 $D=1
M15 GND 612 1343 GND N L=1.8e-07 W=1.17e-06 AD=6.804e-13 AS=4.212e-13 $X=1385500 $Y=940500 $D=1
M16 1344 234 GND GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=6.804e-13 $X=1393500 $Y=942500 $D=1
M17 741 226 1344 GND N L=1.8e-07 W=9.9e-07 AD=5.346e-13 AS=3.564e-13 $X=1399500 $Y=942500 $D=1
M18 1345 818 741 GND N L=1.8e-07 W=9.9e-07 AD=3.564e-13 AS=5.346e-13 $X=1407500 $Y=942500 $D=1
M19 GND 220 1345 GND N L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=3.564e-13 $X=1413500 $Y=942500 $D=1
M20 1346 495 GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.3025e-13 $X=1427500 $Y=1081500 $D=1
M21 1347 111 1346 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=5.508e-13 $X=1433500 $Y=1081500 $D=1
M22 713 20 1347 GND N L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=5.508e-13 $X=1439500 $Y=1081500 $D=1
M23 1348 220 713 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=8.262e-13 $X=1447500 $Y=1081500 $D=1
M24 1349 62 1348 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=5.508e-13 $X=1453500 $Y=1081500 $D=1
M25 GND 34 1349 GND N L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=5.508e-13 $X=1459500 $Y=1081500 $D=1
M26 GND 1337 1336 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.2275e-13 $X=2819500 $Y=40000 $D=1
M27 1350 1339 GND GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=3.078e-13 $X=2827500 $Y=40000 $D=1
M28 1337 1336 1350 GND N L=1.8e-07 W=4.5e-07 AD=7.9785e-13 AS=1.62e-13 $X=2833500 $Y=40000 $D=1
M29 1351 1089 1337 GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.9785e-13 $X=2842000 $Y=29500 $D=1
M30 GND 1338 1351 GND N L=1.8e-07 W=1.53e-06 AD=8.3025e-13 AS=5.508e-13 $X=2848000 $Y=29500 $D=1
M31 GND i_clock 1338 GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=4.9005e-13 $X=2865000 $Y=30500 $D=1
M32 1339 1338 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.994e-13 $X=2873000 $Y=30500 $D=1
M33 1352 1339 GND GND N L=1.8e-07 W=1.53e-06 AD=5.508e-13 AS=7.5735e-13 $X=2889000 $Y=35000 $D=1
M34 1340 1337 1352 GND N L=1.8e-07 W=1.53e-06 AD=7.9785e-13 AS=5.508e-13 $X=2895000 $Y=35000 $D=1
M35 1353 1338 1340 GND N L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=7.9785e-13 $X=2903500 $Y=45000 $D=1
M36 GND 1341 1353 GND N L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=1.62e-13 $X=2909500 $Y=45000 $D=1
M37 1341 1340 GND GND N L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=3.078e-13 $X=2917500 $Y=45000 $D=1
M38 GND 1340 1133 GND N L=1.8e-07 W=9.9e-07 AD=5.994e-13 AS=4.9005e-13 $X=2932500 $Y=26000 $D=1
M39 1114 1133 GND GND N L=1.8e-07 W=9.9e-07 AD=4.9005e-13 AS=5.994e-13 $X=2940500 $Y=26000 $D=1
M40 1354 1299 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.46205e-12 $X=163500 $Y=219500 $D=0
M41 1355 406 1354 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.0368e-12 $X=169500 $Y=219500 $D=0
M42 1356 417 1355 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.0368e-12 $X=175500 $Y=219500 $D=0
M43 404 422 1356 VDD P L=1.8e-07 W=2.88e-06 AD=1.38915e-12 AS=1.0368e-12 $X=181500 $Y=219500 $D=0
M44 1357 535 VDD VDD P L=1.8e-07 W=4.41e-06 AD=1.5876e-12 AS=2.23155e-12 $X=730000 $Y=974500 $D=0
M45 1358 575 1357 VDD P L=1.8e-07 W=4.41e-06 AD=1.5876e-12 AS=1.5876e-12 $X=736000 $Y=974500 $D=0
M46 539 31 1358 VDD P L=1.8e-07 W=4.41e-06 AD=2.47455e-12 AS=1.5876e-12 $X=742000 $Y=974500 $D=0
M47 1359 199 539 VDD P L=1.8e-07 W=3.24e-06 AD=1.1664e-12 AS=2.47455e-12 $X=750500 $Y=987500 $D=0
M48 VDD 194 1359 VDD P L=1.8e-07 W=3.24e-06 AD=1.8225e-12 AS=1.1664e-12 $X=756500 $Y=987500 $D=0
M49 539 584 VDD VDD P L=1.8e-07 W=1.62e-06 AD=7.8975e-13 AS=1.8225e-12 $X=765000 $Y=987500 $D=0
M50 VDD 1331 659 VDD P L=1.8e-07 W=9.9e-07 AD=5.6295e-13 AS=4.9005e-13 $X=963500 $Y=982500 $D=0
M51 1332 224 1331 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=7.5735e-13 $X=979500 $Y=982500 $D=0
M52 VDD 649 1332 VDD P L=1.8e-07 W=1.53e-06 AD=8.91e-13 AS=8.262e-13 $X=987500 $Y=982500 $D=0
M53 1332 205 VDD VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.91e-13 $X=995500 $Y=982500 $D=0
M54 VDD 265 1333 VDD P L=1.8e-07 W=2.34e-06 AD=1.3284e-12 AS=1.12185e-12 $X=1379500 $Y=989500 $D=0
M55 1333 612 VDD VDD P L=1.8e-07 W=2.34e-06 AD=1.215e-12 AS=1.3284e-12 $X=1387500 $Y=989500 $D=0
M56 1334 234 1333 VDD P L=1.8e-07 W=2.07e-06 AD=1.1178e-12 AS=1.215e-12 $X=1395500 $Y=989500 $D=0
M57 1333 226 1334 VDD P L=1.8e-07 W=2.07e-06 AD=1.02465e-12 AS=1.1178e-12 $X=1403500 $Y=989500 $D=0
M58 741 818 1334 VDD P L=1.8e-07 W=2.07e-06 AD=1.1178e-12 AS=1.02465e-12 $X=1419500 $Y=989500 $D=0
M59 1334 220 741 VDD P L=1.8e-07 W=2.07e-06 AD=1.02465e-12 AS=1.1178e-12 $X=1427500 $Y=989500 $D=0
M60 1335 495 VDD VDD P L=1.8e-07 W=1.8e-06 AD=9.72e-13 AS=9.2745e-13 $X=1427500 $Y=1133500 $D=0
M61 VDD 111 1335 VDD P L=1.8e-07 W=1.8e-06 AD=1.0368e-12 AS=9.72e-13 $X=1435500 $Y=1133500 $D=0
M62 1335 20 VDD VDD P L=1.8e-07 W=1.8e-06 AD=9.234e-13 AS=1.0368e-12 $X=1443500 $Y=1133500 $D=0
M63 713 220 1335 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=9.234e-13 $X=1451500 $Y=1133500 $D=0
M64 1335 62 713 VDD P L=1.8e-07 W=1.53e-06 AD=8.262e-13 AS=8.262e-13 $X=1459500 $Y=1133500 $D=0
M65 713 34 1335 VDD P L=1.8e-07 W=1.53e-06 AD=7.5735e-13 AS=8.262e-13 $X=1467500 $Y=1133500 $D=0
M66 VDD 1337 1336 VDD P L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=2.2275e-13 $X=2819500 $Y=73500 $D=0
M67 1360 1338 VDD VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=3.078e-13 $X=2827500 $Y=73500 $D=0
M68 1337 1336 1360 VDD P L=1.8e-07 W=4.5e-07 AD=1.42965e-12 AS=1.62e-13 $X=2833500 $Y=73500 $D=0
M69 1361 1089 1337 VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.42965e-12 $X=2842000 $Y=67500 $D=0
M70 VDD 1339 1361 VDD P L=1.8e-07 W=2.88e-06 AD=1.45395e-12 AS=1.0368e-12 $X=2848000 $Y=67500 $D=0
M71 VDD i_clock 1338 VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=2864000 $Y=77500 $D=0
M72 1339 1338 VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=2872000 $Y=77500 $D=0
M73 1362 1338 VDD VDD P L=1.8e-07 W=2.88e-06 AD=1.0368e-12 AS=1.46205e-12 $X=2888000 $Y=67500 $D=0
M74 1340 1337 1362 VDD P L=1.8e-07 W=2.88e-06 AD=1.42965e-12 AS=1.0368e-12 $X=2894000 $Y=67500 $D=0
M75 1363 1339 1340 VDD P L=1.8e-07 W=4.5e-07 AD=1.62e-13 AS=1.42965e-12 $X=2902500 $Y=82500 $D=0
M76 VDD 1341 1363 VDD P L=1.8e-07 W=4.5e-07 AD=3.078e-13 AS=1.62e-13 $X=2908500 $Y=82500 $D=0
M77 1341 1340 VDD VDD P L=1.8e-07 W=4.5e-07 AD=2.2275e-13 AS=3.078e-13 $X=2916500 $Y=82500 $D=0
M78 VDD 1340 1133 VDD P L=1.8e-07 W=1.98e-06 AD=1.134e-12 AS=9.1935e-13 $X=2932500 $Y=86000 $D=0
M79 1114 1133 VDD VDD P L=1.8e-07 W=1.98e-06 AD=9.1935e-13 AS=1.134e-12 $X=2940500 $Y=86000 $D=0
X80 417 414 437 444 GND VDD mux21 $T=280000 152500 0 0 $X=280000 $Y=152500
X81 427 452 424 423 GND VDD mux21 $T=365500 618500 1 180 $X=312000 $Y=618500
X82 429 427 146 435 GND VDD mux21 $T=328000 783500 0 0 $X=328000 $Y=783500
X83 440 162 448 434 GND VDD mux21 $T=397500 2356500 1 180 $X=344000 $Y=2356500
X84 441 158 449 434 GND VDD mux21 $T=397500 2501500 1 180 $X=344000 $Y=2501500
X85 442 159 450 434 GND VDD mux21 $T=397500 2634500 1 180 $X=344000 $Y=2634500
X86 443 410 459 434 GND VDD mux21 $T=397500 2917500 1 180 $X=344000 $Y=2917500
X87 445 433 453 434 GND VDD mux21 $T=405500 2784500 1 180 $X=352000 $Y=2784500
X88 452 468 154 439 GND VDD mux21 $T=421500 618500 1 180 $X=368000 $Y=618500
X89 458 157 470 125 GND VDD mux21 $T=453500 2223500 1 180 $X=400000 $Y=2223500
X90 448 160 476 i_valid GND VDD mux21 $T=400000 2356500 0 0 $X=400000 $Y=2356500
X91 449 454 219 i_valid GND VDD mux21 $T=400000 2501500 0 0 $X=400000 $Y=2501500
X92 450 455 685 i_valid GND VDD mux21 $T=400000 2634500 0 0 $X=400000 $Y=2634500
X93 459 446 184 i_valid GND VDD mux21 $T=453500 2917500 1 180 $X=400000 $Y=2917500
X94 453 3 568 i_valid GND VDD mux21 $T=408000 2784500 0 0 $X=408000 $Y=2784500
X95 468 497 457 1302 GND VDD mux21 $T=469500 783500 1 180 $X=416000 $Y=783500
X96 460 466 486 8 GND VDD mux21 $T=440000 1474500 0 0 $X=440000 $Y=1474500
X97 470 7 496 i_valid GND VDD mux21 $T=456000 2223500 0 0 $X=456000 $Y=2223500
X98 484 178 170 168 GND VDD mux21 $T=509500 2501500 1 180 $X=456000 $Y=2501500
X99 473 475 173 i_valid GND VDD mux21 $T=464000 2081500 0 0 $X=464000 $Y=2081500
X100 483 166 541 434 GND VDD mux21 $T=464000 2784500 0 0 $X=464000 $Y=2784500
X101 172 481 185 174 GND VDD mux21 $T=525500 783500 1 180 $X=472000 $Y=783500
X102 486 482 182 i_valid GND VDD mux21 $T=549500 1474500 1 180 $X=496000 $Y=1474500
X103 5 14 177 176 GND VDD mux21 $T=573500 461500 1 180 $X=520000 $Y=461500
X104 497 1305 163 485 GND VDD mux21 $T=581500 783500 1 180 $X=528000 $Y=783500
X105 502 41 523 8 GND VDD mux21 $T=613500 7000 1 180 $X=560000 $Y=7000
X106 523 520 193 i_valid GND VDD mux21 $T=669500 7000 1 180 $X=616000 $Y=7000
X107 506 183 533 8 GND VDD mux21 $T=616000 1666500 0 0 $X=616000 $Y=1666500
X108 1305 642 530 190 GND VDD mux21 $T=685500 1200500 1 180 $X=632000 $Y=1200500
X109 514 522 546 187 GND VDD mux21 $T=640000 1057500 0 0 $X=640000 $Y=1057500
X110 533 436 525 i_valid GND VDD mux21 $T=709500 1807500 1 180 $X=656000 $Y=1807500
X111 582 550 1306 534 GND VDD mux21 $T=664000 2501500 0 0 $X=664000 $Y=2501500
X112 412 532 549 176 GND VDD mux21 $T=680000 328500 0 0 $X=680000 $Y=328500
X113 549 109 543 223 GND VDD mux21 $T=749500 152500 1 180 $X=696000 $Y=152500
X114 541 545 639 i_valid GND VDD mux21 $T=712000 2917500 0 0 $X=712000 $Y=2917500
X115 188 i_pixel_bot[15] 76 195 GND VDD mux21 $T=797500 2081500 1 180 $X=744000 $Y=2081500
X116 28 569 198 565 GND VDD mux21 $T=829500 1948500 1 180 $X=776000 $Y=1948500
X117 576 586 592 566 GND VDD mux21 $T=845500 7000 1 180 $X=792000 $Y=7000
X118 610 583 571 573 GND VDD mux21 $T=792000 1341500 0 0 $X=792000 $Y=1341500
X119 583 580 224 588 GND VDD mux21 $T=861500 1200500 1 180 $X=808000 $Y=1200500
X120 198 211 207 613 GND VDD mux21 $T=893500 1807500 1 180 $X=840000 $Y=1807500
X121 503 630 594 634 GND VDD mux21 $T=933500 2917500 1 180 $X=880000 $Y=2917500
X122 608 517 487 223 GND VDD mux21 $T=896000 328500 0 0 $X=896000 $Y=328500
X123 527 47 206 601 GND VDD mux21 $T=981500 2784500 1 180 $X=928000 $Y=2784500
X124 620 628 608 36 GND VDD mux21 $T=997500 461500 1 180 $X=944000 $Y=461500
X125 626 i_pixel_bot[9] 615 623 GND VDD mux21 $T=968000 2223500 0 0 $X=968000 $Y=2223500
X126 631 628 716 648 GND VDD mux21 $T=1045500 328500 1 180 $X=992000 $Y=328500
X127 645 722 627 i_valid GND VDD mux21 $T=1053500 1341500 1 180 $X=1000000 $Y=1341500
X128 553 1310 660 36 GND VDD mux21 $T=1016000 618500 0 0 $X=1016000 $Y=618500
X129 768 i_pixel_bot[17] 652 636 GND VDD mux21 $T=1024000 1807500 0 0 $X=1024000 $Y=1807500
X130 724 i_pixel_top[17] 662 646 GND VDD mux21 $T=1048000 2356500 0 0 $X=1048000 $Y=2356500
X131 225 664 641 21 GND VDD mux21 $T=1101500 2784500 1 180 $X=1048000 $Y=2784500
X132 681 59 645 8 GND VDD mux21 $T=1056000 1341500 0 0 $X=1056000 $Y=1341500
X133 479 643 656 36 GND VDD mux21 $T=1064000 461500 0 0 $X=1064000 $Y=461500
X134 660 221 217 223 GND VDD mux21 $T=1125500 618500 1 180 $X=1072000 $Y=618500
X135 671 39 653 8 GND VDD mux21 $T=1080000 152500 0 0 $X=1080000 $Y=152500
X136 656 101 668 223 GND VDD mux21 $T=1120000 461500 0 0 $X=1120000 $Y=461500
X137 678 673 680 703 GND VDD mux21 $T=1181500 1200500 1 180 $X=1128000 $Y=1200500
X138 252 701 654 26 GND VDD mux21 $T=1205500 2081500 1 180 $X=1152000 $Y=2081500
X139 981 228 687 679 GND VDD mux21 $T=1245500 1474500 1 180 $X=1192000 $Y=1474500
X140 684 689 736 696 GND VDD mux21 $T=1200000 328500 0 0 $X=1200000 $Y=328500
X141 518 233 714 36 GND VDD mux21 $T=1253500 618500 1 180 $X=1200000 $Y=618500
X142 714 136 237 223 GND VDD mux21 $T=1309500 618500 1 180 $X=1256000 $Y=618500
X143 716 33 723 730 GND VDD mux21 $T=1333500 461500 1 180 $X=1280000 $Y=461500
X144 723 233 774 745 GND VDD mux21 $T=1365500 783500 1 180 $X=1312000 $Y=783500
X145 670 740 711 747 GND VDD mux21 $T=1320000 2917500 0 0 $X=1320000 $Y=2917500
X146 725 727 243 767 GND VDD mux21 $T=1360000 2634500 0 0 $X=1360000 $Y=2634500
X147 216 46 49 36 GND VDD mux21 $T=1448000 916500 0 0 $X=1448000 $Y=916500
X148 757 661 780 755 GND VDD mux21 $T=1456000 2501500 0 0 $X=1456000 $Y=2501500
X149 42 771 54 36 GND VDD mux21 $T=1488000 1057500 0 0 $X=1488000 $Y=1057500
X150 775 773 822 795 GND VDD mux21 $T=1573500 461500 1 180 $X=1520000 $Y=461500
X151 941 778 252 803 GND VDD mux21 $T=1560000 2356500 0 0 $X=1560000 $Y=2356500
X152 799 267 806 123 GND VDD mux21 $T=1653500 7000 1 180 $X=1600000 $Y=7000
X153 796 247 855 53 GND VDD mux21 $T=1624000 2917500 0 0 $X=1624000 $Y=2917500
X154 63 820 784 257 GND VDD mux21 $T=1685500 1948500 1 180 $X=1632000 $Y=1948500
X155 801 46 812 51 GND VDD mux21 $T=1640000 916500 0 0 $X=1640000 $Y=916500
X156 806 743 992 i_valid GND VDD mux21 $T=1656000 7000 0 0 $X=1656000 $Y=7000
X157 825 792 i_pixel_top[21] 260 GND VDD mux21 $T=1664000 2784500 0 0 $X=1664000 $Y=2784500
X158 812 818 881 823 GND VDD mux21 $T=1680000 1057500 0 0 $X=1680000 $Y=1057500
X159 54 52 265 809 GND VDD mux21 $T=1696000 916500 0 0 $X=1696000 $Y=916500
X160 603 884 840 294 GND VDD mux21 $T=1789500 1057500 1 180 $X=1736000 $Y=1057500
X161 270 849 817 843 GND VDD mux21 $T=1789500 1807500 1 180 $X=1736000 $Y=1807500
X162 840 111 833 809 GND VDD mux21 $T=1752000 916500 0 0 $X=1752000 $Y=916500
X163 839 876 845 848 GND VDD mux21 $T=1792000 461500 0 0 $X=1792000 $Y=461500
X164 854 841 i_pixel_bot[3] 868 GND VDD mux21 $T=1792000 2634500 0 0 $X=1792000 $Y=2634500
X165 92 850 270 274 GND VDD mux21 $T=1869500 1948500 1 180 $X=1816000 $Y=1948500
X166 874 854 888 859 GND VDD mux21 $T=1840000 2784500 0 0 $X=1840000 $Y=2784500
X167 556 875 886 294 GND VDD mux21 $T=1856000 916500 0 0 $X=1856000 $Y=916500
X168 352 64 872 870 GND VDD mux21 $T=1949500 1666500 1 180 $X=1896000 $Y=1666500
X169 215 874 i_pixel_bot[5] 277 GND VDD mux21 $T=1896000 2784500 0 0 $X=1896000 $Y=2784500
X170 886 917 289 809 GND VDD mux21 $T=1920000 618500 0 0 $X=1920000 $Y=618500
X171 930 65 948 123 GND VDD mux21 $T=1928000 7000 0 0 $X=1928000 $Y=7000
X172 1010 889 1312 883 GND VDD mux21 $T=1981500 1474500 1 180 $X=1928000 $Y=1474500
X173 333 i_pixel_bot[19] 828 69 GND VDD mux21 $T=2005500 1807500 1 180 $X=1952000 $Y=1807500
X174 896 904 895 910 GND VDD mux21 $T=2021500 461500 1 180 $X=1968000 $Y=461500
X175 649 922 903 294 GND VDD mux21 $T=1984000 783500 0 0 $X=1984000 $Y=783500
X176 34 269 931 294 GND VDD mux21 $T=1984000 1057500 0 0 $X=1984000 $Y=1057500
X177 903 956 929 809 GND VDD mux21 $T=2008000 618500 0 0 $X=2008000 $Y=618500
X178 962 869 909 892 GND VDD mux21 $T=2040000 2501500 0 0 $X=2040000 $Y=2501500
X179 906 i_pixel_bot[13] 932 934 GND VDD mux21 $T=2141500 2081500 1 180 $X=2088000 $Y=2081500
X180 918 922 935 928 GND VDD mux21 $T=2104000 916500 0 0 $X=2104000 $Y=916500
X181 940 323 860 i_valid GND VDD mux21 $T=2165500 1666500 1 180 $X=2112000 $Y=1666500
X182 904 929 938 961 GND VDD mux21 $T=2128000 461500 0 0 $X=2128000 $Y=461500
X183 960 942 877 921 GND VDD mux21 $T=2136000 618500 0 0 $X=2136000 $Y=618500
X184 937 312 933 116 GND VDD mux21 $T=2197500 2784500 1 180 $X=2144000 $Y=2784500
X185 959 315 940 129 GND VDD mux21 $T=2221500 1666500 1 180 $X=2168000 $Y=1666500
X186 945 309 947 116 GND VDD mux21 $T=2221500 2634500 1 180 $X=2168000 $Y=2634500
X187 942 317 1106 67 GND VDD mux21 $T=2192000 618500 0 0 $X=2192000 $Y=618500
X188 947 950 974 i_valid GND VDD mux21 $T=2224000 2634500 0 0 $X=2224000 $Y=2634500
X189 963 70 965 972 GND VDD mux21 $T=2309500 328500 1 180 $X=2256000 $Y=328500
X190 1007 91 1029 972 GND VDD mux21 $T=2365500 328500 1 180 $X=2312000 $Y=328500
X191 988 90 990 972 GND VDD mux21 $T=2421500 7000 1 180 $X=2368000 $Y=7000
X192 1005 900 1012 972 GND VDD mux21 $T=2384000 618500 0 0 $X=2384000 $Y=618500
X193 1033 997 94 1002 GND VDD mux21 $T=2469500 2081500 1 180 $X=2416000 $Y=2081500
X194 990 995 332 i_valid GND VDD mux21 $T=2424000 7000 0 0 $X=2424000 $Y=7000
X195 996 74 1014 972 GND VDD mux21 $T=2440000 152500 0 0 $X=2440000 $Y=152500
X196 1000 322 1051 129 GND VDD mux21 $T=2472000 1474500 0 0 $X=2472000 $Y=1474500
X197 1052 326 1069 116 GND VDD mux21 $T=2525500 2917500 1 180 $X=2472000 $Y=2917500
X198 1015 72 1064 972 GND VDD mux21 $T=2496000 152500 0 0 $X=2496000 $Y=152500
X199 1048 339 1006 336 GND VDD mux21 $T=2549500 1200500 1 180 $X=2496000 $Y=1200500
X200 345 99 1016 341 GND VDD mux21 $T=2544000 1948500 0 0 $X=2544000 $Y=1948500
X201 1014 1021 340 i_valid GND VDD mux21 $T=2613500 328500 1 180 $X=2560000 $Y=328500
X202 347 1033 i_pixel_bot[13] 1049 GND VDD mux21 $T=2653500 2081500 1 180 $X=2600000 $Y=2081500
X203 1088 1025 1031 1055 GND VDD mux21 $T=2661500 2356500 1 180 $X=2608000 $Y=2356500
X204 1029 1032 1040 i_valid GND VDD mux21 $T=2616000 328500 0 0 $X=2616000 $Y=328500
X205 1051 955 1222 i_valid GND VDD mux21 $T=2688000 1474500 0 0 $X=2688000 $Y=1474500
X206 1096 352 i_pixel_top[12] 991 GND VDD mux21 $T=2757500 1341500 1 180 $X=2704000 $Y=1341500
X207 1130 1072 346 i_valid GND VDD mux21 $T=2720000 328500 0 0 $X=2720000 $Y=328500
X208 1069 1065 1071 i_valid GND VDD mux21 $T=2773500 2917500 1 180 $X=2720000 $Y=2917500
X209 1064 1068 361 i_valid GND VDD mux21 $T=2744000 152500 0 0 $X=2744000 $Y=152500
X210 1038 1084 1086 1070 GND VDD mux21 $T=2813500 916500 1 180 $X=2760000 $Y=916500
X211 1090 357 310 i_valid GND VDD mux21 $T=2821500 783500 1 180 $X=2768000 $Y=783500
X212 1085 1083 1080 i_valid GND VDD mux21 $T=2837500 2356500 1 180 $X=2784000 $Y=2356500
X213 1132 118 1090 123 GND VDD mux21 $T=2877500 783500 1 180 $X=2824000 $Y=783500
X214 1108 1121 1095 i_valid GND VDD mux21 $T=2893500 2356500 1 180 $X=2840000 $Y=2356500
X215 1316 363 296 i_valid GND VDD mux21 $T=2888000 618500 0 0 $X=2888000 $Y=618500
X216 1156 334 121 328 GND VDD mux21 $T=2941500 2223500 1 180 $X=2888000 $Y=2223500
X217 1158 313 1108 116 GND VDD mux21 $T=2896000 2356500 0 0 $X=2896000 $Y=2356500
X218 119 1149 1112 366 GND VDD mux21 $T=2912000 1807500 0 0 $X=2912000 $Y=1807500
X219 1118 1138 1316 386 GND VDD mux21 $T=2944000 461500 0 0 $X=2944000 $Y=461500
X220 1124 1110 1130 386 GND VDD mux21 $T=2968000 328500 0 0 $X=2968000 $Y=328500
X221 1168 368 i_pixel_top[14] 1128 GND VDD mux21 $T=3029500 1341500 1 180 $X=2976000 $Y=1341500
X222 1153 1155 1170 i_valid GND VDD mux21 $T=3088000 2917500 0 0 $X=3088000 $Y=2917500
X223 1207 1168 1166 1163 GND VDD mux21 $T=3181500 1341500 1 180 $X=3128000 $Y=1341500
X224 1179 372 1157 1171 GND VDD mux21 $T=3181500 1666500 1 180 $X=3128000 $Y=1666500
X225 121 1167 1202 i_valid GND VDD mux21 $T=3136000 2223500 0 0 $X=3136000 $Y=2223500
X226 1227 374 1180 1174 GND VDD mux21 $T=3152000 2917500 0 0 $X=3152000 $Y=2917500
X227 1191 376 132 328 GND VDD mux21 $T=3253500 2356500 1 180 $X=3200000 $Y=2356500
X228 1218 380 1142 127 GND VDD mux21 $T=3224000 1200500 0 0 $X=3224000 $Y=1200500
X229 1204 1189 1188 i_valid GND VDD mux21 $T=3285500 1057500 1 180 $X=3232000 $Y=1057500
X230 1288 383 1218 382 GND VDD mux21 $T=3333500 1200500 1 180 $X=3280000 $Y=1200500
X231 1250 381 1259 129 GND VDD mux21 $T=3341500 1057500 1 180 $X=3288000 $Y=1057500
X232 1197 379 1204 386 GND VDD mux21 $T=3296000 916500 0 0 $X=3296000 $Y=916500
X233 1220 1276 375 i_valid GND VDD mux21 $T=3357500 328500 1 180 $X=3304000 $Y=328500
X234 1217 378 1282 123 GND VDD mux21 $T=3312000 152500 0 0 $X=3312000 $Y=152500
X235 1203 128 1223 129 GND VDD mux21 $T=3312000 1474500 0 0 $X=3312000 $Y=1474500
X236 1226 1209 1290 129 GND VDD mux21 $T=3352000 916500 0 0 $X=3352000 $Y=916500
X237 1228 1268 1220 386 GND VDD mux21 $T=3360000 328500 0 0 $X=3360000 $Y=328500
X238 1244 1229 1317 i_valid GND VDD mux21 $T=3453500 783500 1 180 $X=3400000 $Y=783500
X239 1249 138 1240 1246 GND VDD mux21 $T=3453500 1807500 1 180 $X=3400000 $Y=1807500
X240 1271 1243 1211 1234 GND VDD mux21 $T=3416000 2501500 0 0 $X=3416000 $Y=2501500
X241 132 1239 1264 i_valid GND VDD mux21 $T=3448000 2356500 0 0 $X=3448000 $Y=2356500
X242 1235 393 1244 386 GND VDD mux21 $T=3456000 783500 0 0 $X=3456000 $Y=783500
X243 1318 1248 1252 1254 GND VDD mux21 $T=3488000 2784500 0 0 $X=3488000 $Y=2784500
X244 1259 1255 1283 i_valid GND VDD mux21 $T=3549500 1200500 1 180 $X=3496000 $Y=1200500
X245 1253 1294 1281 386 GND VDD mux21 $T=3512000 783500 0 0 $X=3512000 $Y=783500
X246 1257 1269 1258 1279 GND VDD mux21 $T=3565500 1341500 1 180 $X=3512000 $Y=1341500
X247 1269 1267 399 1273 GND VDD mux21 $T=3552000 1200500 0 0 $X=3552000 $Y=1200500
X248 1281 1296 1277 i_valid GND VDD mux21 $T=3621500 783500 1 180 $X=3568000 $Y=783500
X249 1282 369 401 i_valid GND VDD mux21 $T=3608000 328500 0 0 $X=3608000 $Y=328500
X250 399 1295 1288 1297 GND VDD mux21 $T=3661500 1200500 1 180 $X=3608000 $Y=1200500
X251 1290 1291 1319 i_valid GND VDD mux21 $T=3632000 916500 0 0 $X=3632000 $Y=916500
X252 150 1298 GND VDD inv01 $T=177000 618500 1 180 $X=152000 $Y=618500
X253 436 408 GND VDD inv01 $T=152000 1474500 0 0 $X=152000 $Y=1474500
X254 436 409 GND VDD inv01 $T=152000 1666500 0 0 $X=152000 $Y=1666500
X255 150 407 GND VDD inv01 $T=184000 618500 0 0 $X=184000 $Y=618500
X256 165 415 GND VDD inv01 $T=297000 7000 1 180 $X=272000 $Y=7000
X257 12 419 GND VDD inv01 $T=353000 328500 1 180 $X=328000 $Y=328500
X258 429 426 GND VDD inv01 $T=369000 916500 1 180 $X=344000 $Y=916500
X259 16 457 GND VDD inv01 $T=384000 783500 0 0 $X=384000 $Y=783500
X260 12 169 GND VDD inv01 $T=432000 328500 0 0 $X=432000 $Y=328500
X261 85 434 GND VDD inv01 $T=481000 2356500 1 180 $X=456000 $Y=2356500
X262 171 170 GND VDD inv01 $T=456000 2634500 0 0 $X=456000 $Y=2634500
X263 498 478 GND VDD inv01 $T=537000 1057500 1 180 $X=512000 $Y=1057500
X264 480 515 GND VDD inv01 $T=520000 152500 0 0 $X=520000 $Y=152500
X265 489 218 GND VDD inv01 $T=544000 916500 0 0 $X=544000 $Y=916500
X266 526 499 GND VDD inv01 $T=593000 2081500 1 180 $X=568000 $Y=2081500
X267 551 14 GND VDD inv01 $T=576000 461500 0 0 $X=576000 $Y=461500
X268 436 183 GND VDD inv01 $T=584000 1666500 0 0 $X=584000 $Y=1666500
X269 188 512 GND VDD inv01 $T=657000 2501500 1 180 $X=632000 $Y=2501500
X270 537 513 GND VDD inv01 $T=665000 2784500 1 180 $X=640000 $Y=2784500
X271 32 532 GND VDD inv01 $T=648000 328500 0 0 $X=648000 $Y=328500
X272 153 529 GND VDD inv01 $T=648000 618500 0 0 $X=648000 $Y=618500
X273 i_valid 175 GND VDD inv01 $T=689000 152500 1 180 $X=664000 $Y=152500
X274 125 85 GND VDD inv01 $T=664000 1341500 0 0 $X=664000 $Y=1341500
X275 529 196 GND VDD inv01 $T=680000 618500 0 0 $X=680000 $Y=618500
X276 189 530 GND VDD inv01 $T=713000 1200500 1 180 $X=688000 $Y=1200500
X277 554 191 GND VDD inv01 $T=737000 2081500 1 180 $X=712000 $Y=2081500
X278 577 569 GND VDD inv01 $T=744000 1948500 0 0 $X=744000 $Y=1948500
X279 30 223 GND VDD inv01 $T=752000 152500 0 0 $X=752000 $Y=152500
X280 30 552 GND VDD inv01 $T=777000 618500 1 180 $X=752000 $Y=618500
X281 12 29 GND VDD inv01 $T=825000 783500 1 180 $X=800000 $Y=783500
X282 595 638 GND VDD inv01 $T=832000 783500 0 0 $X=832000 $Y=783500
X283 543 586 GND VDD inv01 $T=873000 7000 1 180 $X=848000 $Y=7000
X284 85 8 GND VDD inv01 $T=848000 1341500 0 0 $X=848000 $Y=1341500
X285 591 776 GND VDD inv01 $T=872000 461500 0 0 $X=872000 $Y=461500
X286 150 15 GND VDD inv01 $T=872000 1057500 0 0 $X=872000 $Y=1057500
X287 776 176 GND VDD inv01 $T=880000 618500 0 0 $X=880000 $Y=618500
X288 218 205 GND VDD inv01 $T=888000 916500 0 0 $X=888000 $Y=916500
X289 208 619 GND VDD inv01 $T=904000 2081500 0 0 $X=904000 $Y=2081500
X290 606 596 GND VDD inv01 $T=937000 1474500 1 180 $X=912000 $Y=1474500
X291 12 20 GND VDD inv01 $T=920000 916500 0 0 $X=920000 $Y=916500
X292 i_pixel_bot[8] 602 GND VDD inv01 $T=961000 2223500 1 180 $X=936000 $Y=2223500
X293 582 641 GND VDD inv01 $T=984000 2784500 0 0 $X=984000 $Y=2784500
X294 1309 621 GND VDD inv01 $T=1017000 783500 1 180 $X=992000 $Y=783500
X295 232 628 GND VDD inv01 $T=1025000 461500 1 180 $X=1000000 $Y=461500
X296 i_pixel_bot[6] 625 GND VDD inv01 $T=1041000 2784500 1 180 $X=1016000 $Y=2784500
X297 254 1310 GND VDD inv01 $T=1049000 783500 1 180 $X=1024000 $Y=783500
X298 33 643 GND VDD inv01 $T=1032000 461500 0 0 $X=1032000 $Y=461500
X299 649 672 GND VDD inv01 $T=1096000 1057500 0 0 $X=1096000 $Y=1057500
X300 666 658 GND VDD inv01 $T=1153000 1474500 1 180 $X=1128000 $Y=1474500
X301 657 675 GND VDD inv01 $T=1128000 1807500 0 0 $X=1128000 $Y=1807500
X302 702 667 GND VDD inv01 $T=1161000 2501500 1 180 $X=1136000 $Y=2501500
X303 674 695 GND VDD inv01 $T=1152000 2223500 0 0 $X=1152000 $Y=2223500
X304 213 687 GND VDD inv01 $T=1160000 1474500 0 0 $X=1160000 $Y=1474500
X305 668 689 GND VDD inv01 $T=1168000 328500 0 0 $X=1168000 $Y=328500
X306 45 150 GND VDD inv01 $T=1193000 618500 1 180 $X=1168000 $Y=618500
X307 i_pixel_bot[16] 688 GND VDD inv01 $T=1168000 1666500 0 0 $X=1168000 $Y=1666500
X308 682 694 GND VDD inv01 $T=1184000 783500 0 0 $X=1184000 $Y=783500
X309 226 680 GND VDD inv01 $T=1209000 1200500 1 180 $X=1184000 $Y=1200500
X310 734 699 GND VDD inv01 $T=1273000 1057500 1 180 $X=1248000 $Y=1057500
X311 241 233 GND VDD inv01 $T=1305000 783500 1 180 $X=1280000 $Y=783500
X312 710 732 GND VDD inv01 $T=1296000 2501500 0 0 $X=1296000 $Y=2501500
X313 34 718 GND VDD inv01 $T=1353000 1057500 1 180 $X=1328000 $Y=1057500
X314 717 235 GND VDD inv01 $T=1361000 1666500 1 180 $X=1336000 $Y=1666500
X315 728 743 GND VDD inv01 $T=1376000 7000 0 0 $X=1376000 $Y=7000
X316 i_pixel_bot[10] 733 GND VDD inv01 $T=1417000 2081500 1 180 $X=1392000 $Y=2081500
X317 743 267 GND VDD inv01 $T=1408000 7000 0 0 $X=1408000 $Y=7000
X318 i_pixel_top[16] 746 GND VDD inv01 $T=1449000 1807500 1 180 $X=1424000 $Y=1807500
X319 i_pixel_top[18] 243 GND VDD inv01 $T=1457000 2356500 1 180 $X=1432000 $Y=2356500
X320 776 36 GND VDD inv01 $T=1481000 461500 1 180 $X=1456000 $Y=461500
X321 217 773 GND VDD inv01 $T=1488000 461500 0 0 $X=1488000 $Y=461500
X322 756 777 GND VDD inv01 $T=1488000 1948500 0 0 $X=1488000 $Y=1948500
X323 248 46 GND VDD inv01 $T=1504000 916500 0 0 $X=1504000 $Y=916500
X324 818 771 GND VDD inv01 $T=1569000 1057500 1 180 $X=1544000 $Y=1057500
X325 776 294 GND VDD inv01 $T=1560000 618500 0 0 $X=1560000 $Y=618500
X326 743 255 GND VDD inv01 $T=1593000 7000 1 180 $X=1568000 $Y=7000
X327 i_pixel_bot[18] 784 GND VDD inv01 $T=1576000 1807500 0 0 $X=1576000 $Y=1807500
X328 i_pixel_top[10] 786 GND VDD inv01 $T=1617000 1474500 1 180 $X=1592000 $Y=1474500
X329 30 809 GND VDD inv01 $T=1640000 618500 0 0 $X=1640000 $Y=618500
X330 809 821 GND VDD inv01 $T=1672000 783500 0 0 $X=1672000 $Y=783500
X331 i_pixel_bot[2] 811 GND VDD inv01 $T=1705000 2356500 1 180 $X=1680000 $Y=2356500
X332 743 846 GND VDD inv01 $T=1712000 152500 0 0 $X=1712000 $Y=152500
X333 826 1311 GND VDD inv01 $T=1777000 1948500 1 180 $X=1752000 $Y=1948500
X334 265 845 GND VDD inv01 $T=1760000 461500 0 0 $X=1760000 $Y=461500
X335 60 850 GND VDD inv01 $T=1784000 1948500 0 0 $X=1784000 $Y=1948500
X336 62 884 GND VDD inv01 $T=1832000 1057500 0 0 $X=1832000 $Y=1057500
X337 908 875 GND VDD inv01 $T=1937000 916500 1 180 $X=1912000 $Y=916500
X338 i_pixel_mid[16] 281 GND VDD inv01 $T=1920000 1807500 0 0 $X=1920000 $Y=1807500
X339 280 o_dir[1] GND VDD inv01 $T=1961000 2917500 1 180 $X=1936000 $Y=2917500
X340 898 1312 GND VDD inv01 $T=1969000 1341500 1 180 $X=1944000 $Y=1341500
X341 i_pixel_bot[4] 888 GND VDD inv01 $T=1977000 2784500 1 180 $X=1952000 $Y=2784500
X342 289 895 GND VDD inv01 $T=2001000 618500 1 180 $X=1976000 $Y=618500
X343 i_pixel_mid[18] 899 GND VDD inv01 $T=2016000 2223500 0 0 $X=2016000 $Y=2223500
X344 300 922 GND VDD inv01 $T=2040000 1057500 0 0 $X=2040000 $Y=1057500
X345 295 902 GND VDD inv01 $T=2065000 1341500 1 180 $X=2040000 $Y=1341500
X346 955 304 GND VDD inv01 $T=2072000 1341500 0 0 $X=2072000 $Y=1341500
X347 936 o_dir[2] GND VDD inv01 $T=2105000 152500 1 180 $X=2080000 $Y=152500
X348 i_pixel_top[22] 923 GND VDD inv01 $T=2112000 2784500 0 0 $X=2112000 $Y=2784500
X349 i_pixel_bot[14] 103 GND VDD inv01 $T=2136000 1807500 0 0 $X=2136000 $Y=1807500
X350 955 830 GND VDD inv01 $T=2193000 1341500 1 180 $X=2168000 $Y=1341500
X351 i_pixel_top[3] 939 GND VDD inv01 $T=2209000 2356500 1 180 $X=2184000 $Y=2356500
X352 i_pixel_top[20] 81 GND VDD inv01 $T=2200000 2784500 0 0 $X=2200000 $Y=2784500
X353 85 116 GND VDD inv01 $T=2216000 2356500 0 0 $X=2216000 $Y=2356500
X354 85 129 GND VDD inv01 $T=2224000 1666500 0 0 $X=2224000 $Y=1666500
X355 i_pixel_bot[19] 949 GND VDD inv01 $T=2257000 2223500 1 180 $X=2232000 $Y=2223500
X356 955 322 GND VDD inv01 $T=2256000 1341500 0 0 $X=2256000 $Y=1341500
X357 85 972 GND VDD inv01 $T=2272000 783500 0 0 $X=2272000 $Y=783500
X358 328 325 GND VDD inv01 $T=2305000 2634500 1 180 $X=2280000 $Y=2634500
X359 85 328 GND VDD inv01 $T=2288000 1057500 0 0 $X=2288000 $Y=1057500
X360 962 979 GND VDD inv01 $T=2369000 2501500 1 180 $X=2344000 $Y=2501500
X361 i_pixel_top[12] 993 GND VDD inv01 $T=2457000 1200500 1 180 $X=2432000 $Y=1200500
X362 i_pixel_top[14] 1006 GND VDD inv01 $T=2464000 1200500 0 0 $X=2464000 $Y=1200500
X363 1010 1315 GND VDD inv01 $T=2553000 1474500 1 180 $X=2528000 $Y=1474500
X364 1045 955 GND VDD inv01 $T=2672000 1341500 0 0 $X=2672000 $Y=1341500
X365 1103 1050 GND VDD inv01 $T=2713000 783500 1 180 $X=2688000 $Y=783500
X366 i_pixel_top[5] 1067 GND VDD inv01 $T=2777000 2501500 1 180 $X=2752000 $Y=2501500
X367 i_pixel_mid[20] 1082 GND VDD inv01 $T=2809000 1948500 1 180 $X=2784000 $Y=1948500
X368 1099 1084 GND VDD inv01 $T=2841000 1057500 1 180 $X=2816000 $Y=1057500
X369 369 1092 GND VDD inv01 $T=2897000 461500 1 180 $X=2872000 $Y=461500
X370 i_pixel_top[13] 1116 GND VDD inv01 $T=2969000 1341500 1 180 $X=2944000 $Y=1341500
X371 i_pixel_bot[21] 1127 GND VDD inv01 $T=2968000 2081500 0 0 $X=2968000 $Y=2081500
X372 367 1141 GND VDD inv01 $T=3065000 916500 1 180 $X=3040000 $Y=916500
X373 1172 386 GND VDD inv01 $T=3072000 916500 0 0 $X=3072000 $Y=916500
X374 1172 123 GND VDD inv01 $T=3176000 783500 0 0 $X=3176000 $Y=783500
X375 i_pixel_mid[22] 1187 GND VDD inv01 $T=3209000 2081500 1 180 $X=3184000 $Y=2081500
X376 125 1172 GND VDD inv01 $T=3225000 1057500 1 180 $X=3200000 $Y=1057500
X377 i_pixel_bot[23] 1180 GND VDD inv01 $T=3233000 2917500 1 180 $X=3208000 $Y=2917500
X378 1237 125 GND VDD inv01 $T=3281000 2223500 1 180 $X=3256000 $Y=2223500
X379 369 124 GND VDD inv01 $T=3297000 328500 1 180 $X=3272000 $Y=328500
X380 369 378 GND VDD inv01 $T=3305000 152500 1 180 $X=3280000 $Y=152500
X381 i_pixel_top[7] 1192 GND VDD inv01 $T=3305000 2501500 1 180 $X=3280000 $Y=2501500
X382 139 1248 GND VDD inv01 $T=3456000 2784500 0 0 $X=3456000 $Y=2784500
X383 392 1267 GND VDD inv01 $T=3464000 1200500 0 0 $X=3464000 $Y=1200500
X384 1245 1243 GND VDD inv01 $T=3497000 2501500 1 180 $X=3472000 $Y=2501500
X385 138 1260 GND VDD inv01 $T=3561000 1666500 1 180 $X=3536000 $Y=1666500
X386 1266 369 GND VDD inv01 $T=3560000 152500 0 0 $X=3560000 $Y=152500
X387 1289 o_dir[0] GND VDD inv01 $T=3624000 783500 0 0 $X=3624000 $Y=783500
X388 400 1285 GND VDD inv01 $T=3649000 2501500 1 180 $X=3624000 $Y=2501500
X389 403 148 146 VDD GND nor02ii $T=193000 783500 1 180 $X=152000 $Y=783500
X390 144 405 403 VDD GND nor02ii $T=193000 916500 1 180 $X=152000 $Y=916500
X391 418 145 144 VDD GND nor02ii $T=193000 1200500 1 180 $X=152000 $Y=1200500
X392 164 413 420 VDD GND nor02ii $T=289000 1666500 1 180 $X=248000 $Y=1666500
X393 431 155 418 VDD GND nor02ii $T=264000 1200500 0 0 $X=264000 $Y=1200500
X394 420 149 467 VDD GND nor02ii $T=321000 1341500 1 180 $X=280000 $Y=1341500
X395 451 432 431 VDD GND nor02ii $T=328000 1341500 0 0 $X=328000 $Y=1341500
X396 429 150 489 VDD GND nor02ii $T=417000 916500 1 180 $X=376000 $Y=916500
X397 467 161 451 VDD GND nor02ii $T=376000 1341500 0 0 $X=376000 $Y=1341500
X398 484 494 1304 VDD GND nor02ii $T=553000 2223500 1 180 $X=512000 $Y=2223500
X399 494 484 519 VDD GND nor02ii $T=561000 2081500 1 180 $X=520000 $Y=2081500
X400 153 176 472 VDD GND nor02ii $T=528000 328500 0 0 $X=528000 $Y=328500
X401 9 183 516 VDD GND nor02ii $T=616000 1341500 0 0 $X=616000 $Y=1341500
X402 205 176 612 VDD GND nor02ii $T=953000 618500 1 180 $X=912000 $Y=618500
X403 i_pixel_bot[8] i_pixel_top[8] 615 VDD GND nor02ii $T=1009000 2501500 1 180 $X=968000 $Y=2501500
X404 677 665 605 VDD GND nor02ii $T=1032000 152500 0 0 $X=1032000 $Y=152500
X405 i_pixel_bot[16] i_pixel_top[0] 652 VDD GND nor02ii $T=1080000 1807500 0 0 $X=1080000 $Y=1807500
X406 i_pixel_top[16] i_pixel_bot[0] 662 VDD GND nor02ii $T=1104000 2356500 0 0 $X=1104000 $Y=2356500
X407 738 700 677 VDD GND nor02ii $T=1136000 152500 0 0 $X=1136000 $Y=152500
X408 242 238 236 VDD GND nor02ii $T=1344000 1200500 0 0 $X=1344000 $Y=1200500
X409 30 104 765 VDD GND nor02ii $T=1472000 618500 0 0 $X=1472000 $Y=618500
X410 794 785 760 VDD GND nor02ii $T=1480000 328500 0 0 $X=1480000 $Y=328500
X411 787 779 772 VDD GND nor02ii $T=1520000 1341500 0 0 $X=1520000 $Y=1341500
X412 761 766 814 VDD GND nor02ii $T=1593000 152500 1 180 $X=1552000 $Y=152500
X413 802 781 787 VDD GND nor02ii $T=1609000 1200500 1 180 $X=1568000 $Y=1200500
X414 807 813 794 VDD GND nor02ii $T=1592000 328500 0 0 $X=1592000 $Y=328500
X415 30 104 283 VDD GND nor02ii $T=1633000 618500 1 180 $X=1592000 $Y=618500
X416 819 815 802 VDD GND nor02ii $T=1616000 1200500 0 0 $X=1616000 $Y=1200500
X417 814 810 807 VDD GND nor02ii $T=1705000 152500 1 180 $X=1664000 $Y=152500
X418 i_pixel_mid[16] i_pixel_mid[0] 816 VDD GND nor02ii $T=1744000 2223500 0 0 $X=1744000 $Y=2223500
X419 858 871 819 VDD GND nor02ii $T=1792000 1200500 0 0 $X=1792000 $Y=1200500
X420 61 846 894 VDD GND nor02ii $T=1849000 152500 1 180 $X=1808000 $Y=152500
X421 269 304 901 VDD GND nor02ii $T=2009000 1200500 1 180 $X=1968000 $Y=1200500
X422 1030 1028 1020 VDD GND nor02ii $T=2560000 618500 0 0 $X=2560000 $Y=618500
X423 1028 1030 999 VDD GND nor02ii $T=2608000 618500 0 0 $X=2608000 $Y=618500
X424 328 i_reset 355 VDD GND nor02ii $T=2761000 783500 1 180 $X=2720000 $Y=783500
X425 98 1092 1074 VDD GND nor02ii $T=2760000 461500 0 0 $X=2760000 $Y=461500
X426 1183 135 1165 VDD GND nor02ii $T=3120000 7000 0 0 $X=3120000 $Y=7000
X427 1169 1162 1176 VDD GND nor02ii $T=3161000 461500 1 180 $X=3120000 $Y=461500
X428 1164 373 1169 VDD GND nor02ii $T=3136000 618500 0 0 $X=3136000 $Y=618500
X429 1176 1181 384 VDD GND nor02ii $T=3273000 461500 1 180 $X=3232000 $Y=461500
X430 384 1242 394 VDD GND nor02ii $T=3497000 461500 1 180 $X=3456000 $Y=461500
X431 1257 1265 1241 VDD GND nor02ii $T=3505000 1474500 1 180 $X=3464000 $Y=1474500
X432 1265 1257 137 VDD GND nor02ii $T=3512000 1474500 0 0 $X=3512000 $Y=1474500
X433 394 1274 134 VDD GND nor02ii $T=3568000 461500 0 0 $X=3568000 $Y=461500
X434 398 1292 396 VDD GND nor02ii $T=3617000 2356500 1 180 $X=3576000 $Y=2356500
X435 1292 398 1286 VDD GND nor02ii $T=3665000 2356500 1 180 $X=3624000 $Y=2356500
X436 408 147 148 GND VDD xnor2 $T=247000 1474500 1 180 $X=184000 $Y=1474500
X437 409 158 149 GND VDD xnor2 $T=247000 1666500 1 180 $X=184000 $Y=1666500
X438 405 144 154 GND VDD xnor2 $T=200000 916500 0 0 $X=200000 $Y=916500
X439 145 418 16 GND VDD xnor2 $T=200000 1200500 0 0 $X=200000 $Y=1200500
X440 409 410 155 GND VDD xnor2 $T=343000 1807500 1 180 $X=280000 $Y=1807500
X441 413 164 209 GND VDD xnor2 $T=359000 1666500 1 180 $X=296000 $Y=1666500
X442 186 165 430 GND VDD xnor2 $T=304000 7000 0 0 $X=304000 $Y=7000
X443 154 425 439 GND VDD xnor2 $T=383000 461500 1 180 $X=320000 $Y=461500
X444 456 437 444 GND VDD xnor2 $T=336000 152500 0 0 $X=336000 $Y=152500
X445 161 467 210 GND VDD xnor2 $T=424000 1341500 0 0 $X=424000 $Y=1341500
X446 563 171 168 GND VDD xnor2 $T=519000 2917500 1 180 $X=456000 $Y=2917500
X447 183 162 504 GND VDD xnor2 $T=543000 1666500 1 180 $X=480000 $Y=1666500
X448 504 511 197 GND VDD xnor2 $T=600000 1474500 0 0 $X=600000 $Y=1474500
X449 519 531 525 GND VDD xnor2 $T=663000 2081500 1 180 $X=600000 $Y=2081500
X450 521 188 531 GND VDD xnor2 $T=640000 2223500 0 0 $X=640000 $Y=2223500
X451 189 538 190 GND VDD xnor2 $T=743000 783500 1 180 $X=680000 $Y=783500
X452 604 546 187 GND VDD xnor2 $T=696000 1057500 0 0 $X=696000 $Y=1057500
X453 551 559 572 GND VDD xnor2 $T=744000 461500 0 0 $X=744000 $Y=461500
X454 76 195 200 GND VDD xnor2 $T=863000 2081500 1 180 $X=800000 $Y=2081500
X455 598 208 577 GND VDD xnor2 $T=895000 1948500 1 180 $X=832000 $Y=1948500
X456 224 614 588 GND VDD xnor2 $T=927000 1200500 1 180 $X=864000 $Y=1200500
X457 616 600 609 GND VDD xnor2 $T=904000 2501500 0 0 $X=904000 $Y=2501500
X458 47 601 630 GND VDD xnor2 $T=999000 2917500 1 180 $X=936000 $Y=2917500
X459 211 613 629 GND VDD xnor2 $T=1007000 1666500 1 180 $X=944000 $Y=1666500
X460 633 654 26 GND VDD xnor2 $T=1063000 2081500 1 180 $X=1000000 $Y=2081500
X461 i_pixel_bot[17] i_pixel_top[1] 636 GND VDD xnor2 $T=1008000 1666500 0 0 $X=1008000 $Y=1666500
X462 666 651 222 GND VDD xnor2 $T=1112000 1341500 0 0 $X=1112000 $Y=1341500
X463 668 101 696 GND VDD xnor2 $T=1176000 461500 0 0 $X=1176000 $Y=461500
X464 770 704 676 GND VDD xnor2 $T=1184000 2917500 0 0 $X=1184000 $Y=2917500
X465 701 26 790 GND VDD xnor2 $T=1271000 2081500 1 180 $X=1208000 $Y=2081500
X466 768 40 555 GND VDD xnor2 $T=1287000 1807500 1 180 $X=1224000 $Y=1807500
X467 742 228 679 GND VDD xnor2 $T=1248000 1474500 0 0 $X=1248000 $Y=1474500
X468 791 706 712 GND VDD xnor2 $T=1256000 1948500 0 0 $X=1256000 $Y=1948500
X469 708 715 721 GND VDD xnor2 $T=1288000 2784500 0 0 $X=1288000 $Y=2784500
X470 724 731 759 GND VDD xnor2 $T=1375000 2356500 1 180 $X=1312000 $Y=2356500
X471 i_pixel_mid[2] i_pixel_bot[1] 710 GND VDD xnor2 $T=1328000 2501500 0 0 $X=1328000 $Y=2501500
X472 241 735 745 GND VDD xnor2 $T=1368000 783500 0 0 $X=1368000 $Y=783500
X473 i_pixel_bot[18] i_pixel_top[2] 40 GND VDD xnor2 $T=1519000 1807500 1 180 $X=1456000 $Y=1807500
X474 766 761 833 GND VDD xnor2 $T=1551000 152500 1 180 $X=1488000 $Y=152500
X475 781 802 248 GND VDD xnor2 $T=1567000 1200500 1 180 $X=1504000 $Y=1200500
X476 785 794 217 GND VDD xnor2 $T=1528000 328500 0 0 $X=1528000 $Y=328500
X477 248 793 51 GND VDD xnor2 $T=1599000 916500 1 180 $X=1536000 $Y=916500
X478 i_pixel_bot[11] i_pixel_top[11] 249 GND VDD xnor2 $T=1607000 2081500 1 180 $X=1544000 $Y=2081500
X479 818 805 823 GND VDD xnor2 $T=1639000 1057500 1 180 $X=1576000 $Y=1057500
X480 810 814 265 GND VDD xnor2 $T=1663000 152500 1 180 $X=1600000 $Y=152500
X481 252 803 869 GND VDD xnor2 $T=1616000 2356500 0 0 $X=1616000 $Y=2356500
X482 816 797 827 GND VDD xnor2 $T=1680000 2223500 0 0 $X=1680000 $Y=2223500
X483 820 257 88 GND VDD xnor2 $T=1688000 1948500 0 0 $X=1688000 $Y=1948500
X484 830 326 779 GND VDD xnor2 $T=1759000 1341500 1 180 $X=1696000 $Y=1341500
X485 255 90 810 GND VDD xnor2 $T=1712000 7000 0 0 $X=1712000 $Y=7000
X486 824 798 861 GND VDD xnor2 $T=1712000 1474500 0 0 $X=1712000 $Y=1474500
X487 846 59 847 GND VDD xnor2 $T=1807000 152500 1 180 $X=1744000 $Y=152500
X488 255 900 785 GND VDD xnor2 $T=2007000 328500 1 180 $X=1944000 $Y=328500
X489 890 894 929 GND VDD xnor2 $T=1952000 152500 0 0 $X=1952000 $Y=152500
X490 64 870 1001 GND VDD xnor2 $T=1952000 1666500 0 0 $X=1952000 $Y=1666500
X491 906 301 266 GND VDD xnor2 $T=2031000 2081500 1 180 $X=1968000 $Y=2081500
X492 898 883 296 GND VDD xnor2 $T=2039000 1341500 1 180 $X=1976000 $Y=1341500
X493 289 915 910 GND VDD xnor2 $T=2024000 461500 0 0 $X=2024000 $Y=461500
X494 300 920 928 GND VDD xnor2 $T=2080000 783500 0 0 $X=2080000 $Y=783500
X495 75 926 958 GND VDD xnor2 $T=2104000 1474500 0 0 $X=2104000 $Y=1474500
X496 830 312 943 GND VDD xnor2 $T=2144000 1200500 0 0 $X=2144000 $Y=1200500
X497 i_pixel_bot[13] i_pixel_top[13] 934 GND VDD xnor2 $T=2231000 1807500 1 180 $X=2168000 $Y=1807500
X498 i_pixel_bot[6] i_pixel_top[22] 966 GND VDD xnor2 $T=2232000 2784500 0 0 $X=2232000 $Y=2784500
X499 322 376 238 GND VDD xnor2 $T=2288000 1341500 0 0 $X=2288000 $Y=1341500
X500 i_pixel_bot[4] i_pixel_top[20] 985 GND VDD xnor2 $T=2312000 2634500 0 0 $X=2312000 $Y=2634500
X501 i_pixel_mid[19] i_pixel_mid[3] 984 GND VDD xnor2 $T=2447000 2223500 1 180 $X=2384000 $Y=2223500
X502 994 1003 1036 GND VDD xnor2 $T=2472000 2784500 0 0 $X=2472000 $Y=2784500
X503 1013 1017 1025 GND VDD xnor2 $T=2567000 2501500 1 180 $X=2504000 $Y=2501500
X504 339 336 1063 GND VDD xnor2 $T=2615000 1200500 1 180 $X=2552000 $Y=1200500
X505 1009 1022 1034 GND VDD xnor2 $T=2560000 1057500 0 0 $X=2560000 $Y=1057500
X506 i_pixel_bot[20] i_pixel_top[4] 1059 GND VDD xnor2 $T=2672000 1807500 0 0 $X=2672000 $Y=1807500
X507 1081 1074 956 GND VDD xnor2 $T=2696000 461500 0 0 $X=2696000 $Y=461500
X508 63 1066 1139 GND VDD xnor2 $T=2720000 1948500 0 0 $X=2720000 $Y=1948500
X509 i_pixel_top[4] i_pixel_top[13] 1091 GND VDD xnor2 $T=2807000 1474500 1 180 $X=2744000 $Y=1474500
X510 354 1099 1070 GND VDD xnor2 $T=2815000 1057500 1 180 $X=2752000 $Y=1057500
X511 1115 1098 917 GND VDD xnor2 $T=2839000 618500 1 180 $X=2776000 $Y=618500
X512 1092 118 1081 GND VDD xnor2 $T=2871000 461500 1 180 $X=2808000 $Y=461500
X513 1136 367 1102 GND VDD xnor2 $T=2943000 783500 1 180 $X=2880000 $Y=783500
X514 124 1138 1115 GND VDD xnor2 $T=3007000 618500 1 180 $X=2944000 $Y=618500
X515 367 1140 1120 GND VDD xnor2 $T=3031000 1057500 1 180 $X=2968000 $Y=1057500
X516 i_pixel_mid[21] i_pixel_bot[22] 1137 GND VDD xnor2 $T=2976000 2634500 0 0 $X=2976000 $Y=2634500
X517 1162 1169 52 GND VDD xnor2 $T=3119000 461500 1 180 $X=3056000 $Y=461500
X518 1149 366 1208 GND VDD xnor2 $T=3064000 1948500 0 0 $X=3064000 $Y=1948500
X519 373 1164 111 GND VDD xnor2 $T=3072000 618500 0 0 $X=3072000 $Y=618500
X520 1152 1150 1184 GND VDD xnor2 $T=3120000 2081500 0 0 $X=3120000 $Y=2081500
X521 1181 1176 106 GND VDD xnor2 $T=3231000 461500 1 180 $X=3168000 $Y=461500
X522 124 379 1181 GND VDD xnor2 $T=3247000 618500 1 180 $X=3184000 $Y=618500
X523 i_pixel_bot[23] 1179 1201 GND VDD xnor2 $T=3247000 1666500 1 180 $X=3184000 $Y=1666500
X524 i_pixel_mid[22] i_pixel_mid[6] 1196 GND VDD xnor2 $T=3192000 2223500 0 0 $X=3192000 $Y=2223500
X525 378 128 371 GND VDD xnor2 $T=3208000 328500 0 0 $X=3208000 $Y=328500
X526 378 381 1182 GND VDD xnor2 $T=3279000 152500 1 180 $X=3216000 $Y=152500
X527 138 1201 1246 GND VDD xnor2 $T=3351000 1666500 1 180 $X=3288000 $Y=1666500
X528 i_pixel_mid[23] 1227 1221 GND VDD xnor2 $T=3359000 2917500 1 180 $X=3296000 $Y=2917500
X529 378 1209 1213 GND VDD xnor2 $T=3312000 618500 0 0 $X=3312000 $Y=618500
X530 i_pixel_top[7] 1207 1232 GND VDD xnor2 $T=3375000 1341500 1 180 $X=3312000 $Y=1341500
X531 1211 1234 1202 GND VDD xnor2 $T=3375000 2501500 1 180 $X=3312000 $Y=2501500
X532 i_pixel_mid[7] 385 1230 GND VDD xnor2 $T=3423000 2634500 1 180 $X=3360000 $Y=2634500
X533 139 1221 390 GND VDD xnor2 $T=3360000 2917500 0 0 $X=3360000 $Y=2917500
X534 1242 384 221 GND VDD xnor2 $T=3392000 461500 0 0 $X=3392000 $Y=461500
X535 1230 1245 1234 GND VDD xnor2 $T=3424000 2634500 0 0 $X=3424000 $Y=2634500
X536 124 393 1242 GND VDD xnor2 $T=3432000 618500 0 0 $X=3432000 $Y=618500
X537 139 1247 1254 GND VDD xnor2 $T=3464000 2917500 0 0 $X=3464000 $Y=2917500
X538 1274 394 136 GND VDD xnor2 $T=3504000 461500 0 0 $X=3504000 $Y=461500
X539 1271 1280 1264 GND VDD xnor2 $T=3504000 2356500 0 0 $X=3504000 $Y=2356500
X540 396 397 1222 GND VDD xnor2 $T=3528000 2223500 0 0 $X=3528000 $Y=2223500
X541 1261 139 397 GND VDD xnor2 $T=3528000 2634500 0 0 $X=3528000 $Y=2634500
X542 1252 1254 400 GND VDD xnor2 $T=3544000 2784500 0 0 $X=3544000 $Y=2784500
X543 399 1273 1319 GND VDD xnor2 $T=3608000 1057500 0 0 $X=3608000 $Y=1057500
X544 1278 138 1320 GND VDD xnor2 $T=3608000 1666500 0 0 $X=3608000 $Y=1666500
X545 124 1294 1274 GND VDD xnor2 $T=3616000 461500 0 0 $X=3616000 $Y=461500
X546 137 1320 401 GND VDD xnor2 $T=3624000 1474500 0 0 $X=3624000 $Y=1474500
X547 5 407 416 GND VDD nand02 $T=200000 461500 0 0 $X=200000 $Y=461500
X548 412 407 1301 GND VDD nand02 $T=273000 461500 1 180 $X=240000 $Y=461500
X549 429 150 421 GND VDD nand02 $T=297000 916500 1 180 $X=264000 $Y=916500
X550 620 407 425 GND VDD nand02 $T=280000 461500 0 0 $X=280000 $Y=461500
X551 421 426 12 GND VDD nand02 $T=304000 916500 0 0 $X=304000 $Y=916500
X552 479 407 1303 GND VDD nand02 $T=473000 461500 1 180 $X=440000 $Y=461500
X553 183 493 180 GND VDD nand02 $T=544000 1666500 0 0 $X=544000 $Y=1666500
X554 518 407 490 GND VDD nand02 $T=585000 618500 1 180 $X=552000 $Y=618500
X555 521 188 494 GND VDD nand02 $T=593000 2223500 1 180 $X=560000 $Y=2223500
X556 188 179 521 GND VDD nand02 $T=633000 2223500 1 180 $X=600000 $Y=2223500
X557 526 i_valid 528 GND VDD nand02 $T=689000 1948500 1 180 $X=656000 $Y=1948500
X558 194 199 524 GND VDD nand02 $T=705000 916500 1 180 $X=672000 $Y=916500
X559 553 407 538 GND VDD nand02 $T=745000 618500 1 180 $X=712000 $Y=618500
X560 556 15 1308 GND VDD nand02 $T=753000 1200500 1 180 $X=720000 $Y=1200500
X561 i_pixel_top[16] i_pixel_mid[17] 579 GND VDD nand02 $T=752000 2356500 0 0 $X=752000 $Y=2356500
X562 558 i_pixel_top[23] 563 GND VDD nand02 $T=768000 2917500 0 0 $X=768000 $Y=2917500
X563 589 i_pixel_bot[7] 567 GND VDD nand02 $T=833000 2634500 1 180 $X=800000 $Y=2634500
X564 27 587 584 GND VDD nand02 $T=881000 916500 1 180 $X=848000 $Y=916500
X565 602 i_pixel_top[8] 585 GND VDD nand02 $T=881000 2223500 1 180 $X=848000 $Y=2223500
X566 i_pixel_top[8] i_pixel_top[17] 593 GND VDD nand02 $T=889000 1666500 1 180 $X=856000 $Y=1666500
X567 i_pixel_bot[8] i_pixel_bot[1] 598 GND VDD nand02 $T=897000 2081500 1 180 $X=864000 $Y=2081500
X568 15 603 599 GND VDD nand02 $T=961000 1200500 1 180 $X=928000 $Y=1200500
X569 649 15 614 GND VDD nand02 $T=1001000 1200500 1 180 $X=968000 $Y=1200500
X570 216 15 632 GND VDD nand02 $T=1016000 1057500 0 0 $X=1016000 $Y=1057500
X571 42 15 697 GND VDD nand02 $T=1056000 1057500 0 0 $X=1056000 $Y=1057500
X572 i_pixel_bot[17] i_pixel_mid[16] 663 GND VDD nand02 $T=1097000 2081500 1 180 $X=1064000 $Y=2081500
X573 i_pixel_top[0] 688 691 GND VDD nand02 $T=1200000 1666500 0 0 $X=1200000 $Y=1666500
X574 i_pixel_bot[0] i_pixel_mid[1] 692 GND VDD nand02 $T=1200000 2634500 0 0 $X=1200000 $Y=2634500
X575 i_pixel_bot[16] i_pixel_bot[9] 764 GND VDD nand02 $T=1320000 1948500 0 0 $X=1320000 $Y=1948500
X576 666 i_valid 244 GND VDD nand02 $T=1368000 1341500 0 0 $X=1368000 $Y=1341500
X577 i_pixel_bot[0] 746 729 GND VDD nand02 $T=1417000 1807500 1 180 $X=1384000 $Y=1807500
X578 294 765 45 GND VDD nand02 $T=1553000 618500 1 180 $X=1520000 $Y=618500
X579 i_pixel_top[9] i_pixel_top[0] 824 GND VDD nand02 $T=1624000 1474500 0 0 $X=1624000 $Y=1474500
X580 104 52 838 GND VDD nand02 $T=1720000 618500 0 0 $X=1720000 $Y=618500
X581 826 i_valid 837 GND VDD nand02 $T=1728000 1666500 0 0 $X=1728000 $Y=1666500
X582 i_pixel_top[1] i_pixel_mid[0] 844 GND VDD nand02 $T=1792000 2223500 0 0 $X=1792000 $Y=2223500
X583 267 864 853 GND VDD nand02 $T=1832000 7000 0 0 $X=1832000 $Y=7000
X584 104 111 863 GND VDD nand02 $T=1913000 618500 1 180 $X=1880000 $Y=618500
X585 i_pixel_mid[0] 281 879 GND VDD nand02 $T=1953000 1948500 1 180 $X=1920000 $Y=1948500
X586 104 917 915 GND VDD nand02 $T=2121000 461500 1 180 $X=2088000 $Y=461500
X587 295 i_valid 318 GND VDD nand02 $T=2200000 1057500 0 0 $X=2200000 $Y=1057500
X588 322 1314 317 GND VDD nand02 $T=2241000 1200500 1 180 $X=2208000 $Y=1200500
X589 1048 i_pixel_top[15] 1046 GND VDD nand02 $T=2616000 1200500 0 0 $X=2616000 $Y=1200500
X590 378 1134 1106 GND VDD nand02 $T=2937000 461500 1 180 $X=2904000 $Y=461500
X591 1136 367 1028 GND VDD nand02 $T=2977000 783500 1 180 $X=2944000 $Y=783500
X592 1144 1148 344 GND VDD nand02 $T=2993000 7000 1 180 $X=2960000 $Y=7000
X593 367 1135 1136 GND VDD nand02 $T=3000000 916500 0 0 $X=3000000 $Y=916500
X594 348 i_pixel_bot[15] 1140 GND VDD nand02 $T=3065000 1057500 1 180 $X=3032000 $Y=1057500
X595 1179 i_pixel_bot[23] 1219 GND VDD nand02 $T=3248000 1666500 0 0 $X=3248000 $Y=1666500
X596 1207 i_pixel_top[7] 1236 GND VDD nand02 $T=3376000 1341500 0 0 $X=3376000 $Y=1341500
X597 385 i_pixel_mid[7] 1263 GND VDD nand02 $T=3409000 2501500 1 180 $X=3376000 $Y=2501500
X598 1227 i_pixel_mid[23] 1247 GND VDD nand02 $T=3424000 2917500 0 0 $X=3424000 $Y=2917500
X599 139 1318 1261 GND VDD nand02 $T=3521000 2634500 1 180 $X=3488000 $Y=2634500
X600 1278 138 1265 GND VDD nand02 $T=3593000 1474500 1 180 $X=3560000 $Y=1474500
X601 138 1270 1278 GND VDD nand02 $T=3568000 1666500 0 0 $X=3568000 $Y=1666500
X602 1261 139 398 GND VDD nand02 $T=3625000 2634500 1 180 $X=3592000 $Y=2634500
X603 488 519 175 1304 GND VDD nor03 $T=553000 1948500 1 180 $X=512000 $Y=1948500
X604 511 495 482 183 GND VDD nor03 $T=552000 1474500 0 0 $X=552000 $Y=1474500
X605 544 191 i_pixel_mid[16] 547 GND VDD nor03 $T=696000 1948500 0 0 $X=696000 $Y=1948500
X606 240 235 i_pixel_top[16] 719 GND VDD nor03 $T=1360000 1474500 0 0 $X=1360000 $Y=1474500
X607 834 758 i_pixel_top[0] 750 GND VDD nor03 $T=1520000 1666500 0 0 $X=1520000 $Y=1666500
X608 851 261 263 267 GND VDD nor03 $T=1809000 328500 1 180 $X=1768000 $Y=328500
X609 307 911 i_pixel_top[8] 916 GND VDD nor03 $T=2064000 1666500 0 0 $X=2064000 $Y=1666500
X610 952 320 323 322 GND VDD nor03 $T=2240000 1057500 0 0 $X=2240000 $Y=1057500
X611 327 999 175 1020 GND VDD nor03 $T=2377000 618500 1 180 $X=2336000 $Y=618500
X612 1027 101 221 136 GND VDD nor03 $T=2585000 461500 1 180 $X=2544000 $Y=461500
X613 1044 106 917 52 GND VDD nor03 $T=2689000 461500 1 180 $X=2648000 $Y=461500
X614 1056 107 517 109 GND VDD nor03 $T=2713000 328500 1 180 $X=2672000 $Y=328500
X615 1060 357 111 319 GND VDD nor03 $T=2728000 618500 0 0 $X=2728000 $Y=618500
X616 1098 319 357 378 GND VDD nor03 $T=2881000 618500 1 180 $X=2840000 $Y=618500
X617 1233 137 395 1241 GND VDD nor03 $T=3457000 1474500 1 180 $X=3416000 $Y=1474500
X618 1284 396 395 1286 GND VDD nor03 $T=3633000 2223500 1 180 $X=3592000 $Y=2223500
X619 1298 5 146 1300 VDD GND aoi21 $T=152000 461500 0 0 $X=152000 $Y=461500
X620 156 175 488 469 VDD GND aoi21 $T=464000 1948500 0 0 $X=464000 $Y=1948500
X621 585 597 i_pixel_mid[0] 547 VDD GND aoi21 $T=704000 2223500 0 0 $X=704000 $Y=2223500
X622 15 34 9 580 VDD GND aoi21 $T=801000 1200500 1 180 $X=760000 $Y=1200500
X623 691 655 i_pixel_bot[0] 719 VDD GND aoi21 $T=1329000 1666500 1 180 $X=1288000 $Y=1666500
X624 729 720 i_pixel_bot[16] 750 VDD GND aoi21 $T=1465000 1666500 1 180 $X=1424000 $Y=1666500
X625 879 288 i_pixel_bot[8] 916 VDD GND aoi21 $T=2008000 1948500 0 0 $X=2008000 $Y=1948500
X626 104 319 61 938 VDD GND aoi21 $T=2225000 461500 1 180 $X=2184000 $Y=461500
X627 944 175 327 948 VDD GND aoi21 $T=2200000 152500 0 0 $X=2200000 $Y=152500
X628 135 1183 1133 1216 VDD GND aoi21 $T=3209000 7000 1 180 $X=3168000 $Y=7000
X629 1215 395 1233 1223 VDD GND aoi21 $T=3368000 1474500 0 0 $X=3368000 $Y=1474500
X630 1275 395 1284 388 VDD GND aoi21 $T=3584000 2081500 0 0 $X=3584000 $Y=2081500
X631 148 403 152 146 416 435 GND VDD ICV_1 $T=200000 783500 0 0 $X=200000 $Y=783500
X632 155 431 163 432 451 189 GND VDD ICV_1 $T=312000 1200500 0 0 $X=312000 $Y=1200500
X633 611 207 613 652 636 611 GND VDD ICV_1 $T=896000 1807500 0 0 $X=896000 $Y=1807500
X634 615 623 616 662 646 633 GND VDD ICV_1 $T=920000 2356500 0 0 $X=920000 $Y=2356500
X635 229 702 690 692 710 702 GND VDD ICV_1 $T=1168000 2501500 0 0 $X=1168000 $Y=2501500
X636 i_pixel_mid[22] i_pixel_top[21] 260 i_pixel_mid[20] i_pixel_top[19] 245 GND VDD ICV_1 $T=1664000 2634500 0 0 $X=1664000 $Y=2634500
X637 262 855 53 266 835 789 GND VDD ICV_1 $T=1680000 2917500 0 0 $X=1680000 $Y=2917500
X638 826 264 860 i_pixel_top[2] i_pixel_top[11] 870 GND VDD ICV_1 $T=1768000 1666500 0 0 $X=1768000 $Y=1666500
X639 854 859 855 874 277 835 GND VDD ICV_1 $T=1808000 2917500 0 0 $X=1808000 $Y=2917500
X640 941 953 973 962 969 974 GND VDD ICV_1 $T=2216000 2501500 0 0 $X=2216000 $Y=2501500
X641 80 980 970 989 957 980 GND VDD ICV_1 $T=2232000 1807500 0 0 $X=2232000 $Y=1807500
X642 981 964 332 322 334 752 GND VDD ICV_1 $T=2344000 1474500 0 0 $X=2344000 $Y=1474500
X643 92 998 335 99 341 338 GND VDD ICV_1 $T=2416000 1948500 0 0 $X=2416000 $Y=1948500
X644 1010 1023 346 347 1039 351 GND VDD ICV_1 $T=2560000 1474500 0 0 $X=2560000 $Y=1474500
X645 1033 1049 356 i_pixel_mid[20] i_pixel_mid[4] 1075 GND VDD ICV_1 $T=2656000 2081500 0 0 $X=2656000 $Y=2081500
X646 1079 1075 1109 i_pixel_mid[20] i_pixel_bot[21] 364 GND VDD ICV_1 $T=2840000 2081500 0 0 $X=2840000 $Y=2081500
X647 367 1175 1117 i_pixel_bot[15] 348 1175 GND VDD ICV_1 $T=3072000 1057500 0 0 $X=3072000 $Y=1057500
X648 124 1110 373 124 1268 1162 GND VDD ICV_1 $T=3080000 328500 0 0 $X=3080000 $Y=328500
X649 1269 1279 1283 140 1295 1297 GND VDD ICV_1 $T=3568000 1341500 0 0 $X=3568000 $Y=1341500
X650 1272 1262 1287 1293 1287 1295 GND VDD ICV_1 $T=3576000 1807500 0 0 $X=3576000 $Y=1807500
X651 414 444 406 VDD GND xor2 $T=279000 152500 1 180 $X=208000 $Y=152500
X652 481 174 474 VDD GND xor2 $T=543000 916500 1 180 $X=472000 $Y=916500
X653 594 634 184 VDD GND xor2 $T=879000 2917500 1 180 $X=808000 $Y=2917500
X654 711 747 685 VDD GND xor2 $T=1319000 2917500 1 180 $X=1248000 $Y=2917500
X655 921 67 306 VDD GND xor2 $T=2135000 618500 1 180 $X=2064000 $Y=618500
X656 329 975 971 VDD GND xor2 $T=2375000 783500 1 180 $X=2304000 $Y=783500
X657 353 350 1040 VDD GND xor2 $T=2727000 618500 1 180 $X=2656000 $Y=618500
X658 1088 359 1095 VDD GND xor2 $T=2855000 2501500 1 180 $X=2784000 $Y=2501500
X659 1142 127 1188 VDD GND xor2 $T=3223000 1200500 1 180 $X=3152000 $Y=1200500
X660 1206 1186 1170 VDD GND xor2 $T=3239000 2634500 1 180 $X=3168000 $Y=2634500
X661 1288 1297 1277 VDD GND xor2 $T=3607000 1057500 1 180 $X=3536000 $Y=1057500
X662 414 172 415 430 172 430 1299 GND VDD ICV_2 $T=215000 7000 1 180 $X=152000 $Y=7000
X663 492 192 499 181 492 534 476 GND VDD ICV_2 $T=551000 2356500 1 180 $X=488000 $Y=2356500
X664 673 610 209 618 209 599 618 GND VDD ICV_2 $T=943000 1341500 1 180 $X=880000 $Y=1341500
X665 642 678 210 650 210 632 650 GND VDD ICV_2 $T=1071000 1200500 1 180 $X=1008000 $Y=1200500
X666 749 725 i_pixel_top[19] 245 725 245 708 GND VDD ICV_2 $T=1303000 2634500 1 180 $X=1240000 $Y=2634500
X667 247 757 788 783 757 783 715 GND VDD ICV_2 $T=1479000 2634500 1 180 $X=1416000 $Y=2634500
X668 47 796 835 789 796 789 704 GND VDD ICV_2 $T=1567000 2917500 1 180 $X=1504000 $Y=2917500
X669 876 896 833 885 833 863 885 GND VDD ICV_2 $T=1911000 461500 1 180 $X=1848000 $Y=461500
X670 348 347 103 1039 1054 1016 341 GND VDD ICV_2 $T=2615000 1807500 1 180 $X=2552000 $Y=1807500
X671 1030 1038 1050 349 1038 349 340 GND VDD ICV_2 $T=2631000 783500 1 180 $X=2568000 $Y=783500
X672 1101 1053 1057 1035 1053 1035 1087 GND VDD ICV_2 $T=2679000 2634500 1 180 $X=2616000 $Y=2634500
X673 1146 331 1153 116 1129 1125 1071 GND VDD ICV_2 $T=2839000 2917500 1 180 $X=2776000 $Y=2917500
X674 374 1111 i_pixel_bot[22] 1137 1111 1137 1097 GND VDD ICV_2 $T=2919000 2634500 1 180 $X=2856000 $Y=2634500
X675 1211 1205 1206 1186 1193 1205 1186 GND VDD ICV_2 $T=3303000 2634500 1 180 $X=3240000 $Y=2634500
X676 1292 1271 1285 1280 1263 400 1280 GND VDD ICV_2 $T=3567000 2501500 1 180 $X=3504000 $Y=2501500
X677 539 522 622 498 471 GND VDD ICV_3 $T=544000 1057500 0 0 $X=544000 $Y=1057500
X678 510 436 526 181 182 GND VDD ICV_3 $T=560000 1948500 0 0 $X=560000 $Y=1948500
X679 524 535 539 187 509 GND VDD ICV_3 $T=576000 916500 0 0 $X=576000 $Y=916500
X680 218 153 560 185 174 GND VDD ICV_3 $T=584000 783500 0 0 $X=584000 $Y=783500
X681 492 1306 542 192 181 GND VDD ICV_3 $T=608000 2356500 0 0 $X=608000 $Y=2356500
X682 798 808 i_pixel_top[1] i_pixel_top[10] 798 GND VDD ICV_3 $T=1568000 1666500 0 0 $X=1568000 $Y=1666500
X683 o_edge 324 255 39 890 GND VDD ICV_3 $T=1856000 152500 0 0 $X=1856000 $Y=152500
X684 i_pixel_bot[12] 94 i_pixel_bot[12] i_pixel_top[12] 87 GND VDD ICV_3 $T=2320000 2081500 0 0 $X=2320000 $Y=2081500
X685 i_pixel_bot[20] 1112 1107 356 1078 GND VDD ICV_3 $T=2752000 1666500 0 0 $X=2752000 $Y=1666500
X686 i_pixel_top[15] 1166 368 1128 1194 GND VDD ICV_3 $T=3032000 1341500 0 0 $X=3032000 $Y=1341500
X687 i_pixel_bot[22] 1157 i_pixel_bot[22] i_pixel_top[6] 1151 GND VDD ICV_3 $T=3032000 1666500 0 0 $X=3032000 $Y=1666500
X688 i_valid 395 1238 1256 1272 GND VDD ICV_3 $T=3496000 1948500 0 0 $X=3496000 $Y=1948500
X689 438 i_reset i_clock 1321 o_mode[1] GND VDD dffr $T=337000 1057500 1 180 $X=152000 $Y=1057500
X690 465 i_reset i_clock 147 156 GND VDD dffr $T=337000 1948500 1 180 $X=152000 $Y=1948500
X691 464 i_reset i_clock 151 475 GND VDD dffr $T=337000 2081500 1 180 $X=152000 $Y=2081500
X692 458 i_reset i_clock 157 7 GND VDD dffr $T=337000 2223500 1 180 $X=152000 $Y=2223500
X693 440 i_reset i_clock 162 160 GND VDD dffr $T=337000 2356500 1 180 $X=152000 $Y=2356500
X694 441 i_reset i_clock 158 454 GND VDD dffr $T=337000 2501500 1 180 $X=152000 $Y=2501500
X695 442 i_reset i_clock 159 455 GND VDD dffr $T=337000 2634500 1 180 $X=152000 $Y=2634500
X696 443 i_reset i_clock 410 446 GND VDD dffr $T=337000 2917500 1 180 $X=152000 $Y=2917500
X697 445 i_reset i_clock 433 3 GND VDD dffr $T=345000 2784500 1 180 $X=160000 $Y=2784500
X698 460 i_reset i_clock 466 482 GND VDD dffr $T=248000 1474500 0 0 $X=248000 $Y=1474500
X699 502 i_reset i_clock 41 520 GND VDD dffr $T=553000 7000 1 180 $X=368000 $Y=7000
X700 540 i_reset i_clock 9 495 GND VDD dffr $T=625000 1200500 1 180 $X=440000 $Y=1200500
X701 506 i_reset i_clock 510 1322 GND VDD dffr $T=464000 1807500 0 0 $X=464000 $Y=1807500
X702 483 i_reset i_clock 166 545 GND VDD dffr $T=520000 2917500 0 0 $X=520000 $Y=2917500
X703 671 i_reset i_clock 39 263 GND VDD dffr $T=1177000 7000 1 180 $X=992000 $Y=7000
X704 681 i_reset i_clock 59 722 GND VDD dffr $T=1176000 1341500 0 0 $X=1176000 $Y=1341500
X705 799 i_reset i_clock 728 1323 GND VDD dffr $T=1369000 7000 1 180 $X=1184000 $Y=7000
X706 856 i_reset i_clock 61 261 GND VDD dffr $T=1889000 783500 1 180 $X=1704000 $Y=783500
X707 945 i_reset i_clock 309 950 GND VDD dffr $T=2161000 2634500 1 180 $X=1976000 $Y=2634500
X708 930 i_reset i_clock 65 944 GND VDD dffr $T=2169000 7000 1 180 $X=1984000 $Y=7000
X709 963 i_reset i_clock 70 968 GND VDD dffr $T=2249000 328500 1 180 $X=2064000 $Y=328500
X710 937 i_reset i_clock 312 924 GND VDD dffr $T=2088000 2917500 0 0 $X=2088000 $Y=2917500
X711 988 i_reset i_clock 90 995 GND VDD dffr $T=2176000 7000 0 0 $X=2176000 $Y=7000
X712 996 i_reset i_clock 74 1021 GND VDD dffr $T=2248000 152500 0 0 $X=2248000 $Y=152500
X713 959 i_reset i_clock 315 323 GND VDD dffr $T=2256000 1666500 0 0 $X=2256000 $Y=1666500
X714 325 i_reset i_clock 1324 o_valid GND VDD dffr $T=2280000 2917500 0 0 $X=2280000 $Y=2917500
X715 978 i_reset i_clock 269 320 GND VDD dffr $T=2328000 916500 0 0 $X=2328000 $Y=916500
X716 1005 i_reset i_clock 900 1008 GND VDD dffr $T=2537000 461500 1 180 $X=2352000 $Y=461500
X717 1007 i_reset i_clock 91 1032 GND VDD dffr $T=2553000 328500 1 180 $X=2368000 $Y=328500
X718 986 i_reset i_clock 98 319 GND VDD dffr $T=2376000 783500 0 0 $X=2376000 $Y=783500
X719 1000 i_reset i_clock 1045 1325 GND VDD dffr $T=2480000 1341500 0 0 $X=2480000 $Y=1341500
X720 1052 i_reset i_clock 326 1065 GND VDD dffr $T=2713000 2917500 1 180 $X=2528000 $Y=2917500
X721 1015 i_reset i_clock 72 1068 GND VDD dffr $T=2552000 152500 0 0 $X=2552000 $Y=152500
X722 1094 i_reset i_clock 311 1083 GND VDD dffr $T=2881000 2223500 1 180 $X=2696000 $Y=2223500
X723 1124 i_reset i_clock 1110 1072 GND VDD dffr $T=2961000 328500 1 180 $X=2776000 $Y=328500
X724 1146 i_reset i_clock 331 1155 GND VDD dffr $T=3081000 2917500 1 180 $X=2896000 $Y=2917500
X725 1118 i_reset i_clock 1138 363 GND VDD dffr $T=2912000 152500 0 0 $X=2912000 $Y=152500
X726 1156 i_reset i_clock 334 1167 GND VDD dffr $T=3129000 2223500 1 180 $X=2944000 $Y=2223500
X727 1158 i_reset i_clock 313 1121 GND VDD dffr $T=3137000 2356500 1 180 $X=2952000 $Y=2356500
X728 1132 i_reset i_clock 118 357 GND VDD dffr $T=2984000 783500 0 0 $X=2984000 $Y=783500
X729 1197 i_reset i_clock 379 1189 GND VDD dffr $T=3289000 916500 1 180 $X=3104000 $Y=916500
X730 1203 i_reset i_clock 128 1215 GND VDD dffr $T=3305000 1474500 1 180 $X=3120000 $Y=1474500
X731 1235 i_reset i_clock 393 1229 GND VDD dffr $T=3393000 783500 1 180 $X=3208000 $Y=783500
X732 1216 i_reset i_clock 1183 1326 GND VDD dffr $T=3401000 7000 1 180 $X=3216000 $Y=7000
X733 1191 i_reset i_clock 376 1239 GND VDD dffr $T=3256000 2356500 0 0 $X=3256000 $Y=2356500
X734 1251 i_reset i_clock 1327 1237 GND VDD dffr $T=3288000 2223500 0 0 $X=3288000 $Y=2223500
X735 1250 i_reset i_clock 381 1255 GND VDD dffr $T=3529000 1057500 1 180 $X=3344000 $Y=1057500
X736 1217 i_reset i_clock 1266 1328 GND VDD dffr $T=3368000 152500 0 0 $X=3368000 $Y=152500
X737 1224 i_reset i_clock 314 1275 GND VDD dffr $T=3392000 2081500 0 0 $X=3392000 $Y=2081500
X738 1226 i_reset i_clock 1209 1291 GND VDD dffr $T=3408000 916500 0 0 $X=3408000 $Y=916500
X739 1228 i_reset i_clock 1268 1276 GND VDD dffr $T=3416000 328500 0 0 $X=3416000 $Y=328500
X740 1253 i_reset i_clock 1294 1296 GND VDD dffr $T=3496000 618500 0 0 $X=3496000 $Y=618500
X741 12 294 67 GND VDD and02 $T=1849500 916500 1 180 $X=1808000 $Y=916500
X742 i_valid 328 1251 GND VDD and02 $T=3480000 2223500 0 0 $X=3480000 $Y=2223500
X743 464 151 473 125 409 166 432 GND VDD ICV_4 $T=344000 2081500 0 0 $X=344000 $Y=2081500
X744 49 106 239 223 237 136 748 GND VDD ICV_4 $T=1352000 618500 0 0 $X=1352000 $Y=618500
X745 887 i_pixel_bot[11] 769 249 i_pixel_bot[3] i_pixel_bot[10] 753 GND VDD ICV_4 $T=1424000 2081500 0 0 $X=1424000 $Y=2081500
X746 877 180 853 67 265 838 848 GND VDD ICV_4 $T=1760000 618500 0 0 $X=1760000 $Y=618500
X747 933 924 298 i_valid i_pixel_mid[6] i_pixel_bot[5] 277 GND VDD ICV_4 $T=1968000 2917500 0 0 $X=1968000 $Y=2917500
X748 997 84 i_pixel_bot[11] 316 932 934 262 GND VDD ICV_4 $T=2144000 2081500 0 0 $X=2144000 $Y=2081500
X749 982 i_pixel_top[21] 994 1003 982 966 114 GND VDD ICV_4 $T=2352000 2784500 0 0 $X=2352000 $Y=2784500
X750 1094 311 1085 116 1031 1055 1080 GND VDD ICV_4 $T=2664000 2356500 0 0 $X=2664000 $Y=2356500
X751 1206 1145 1129 1125 1101 1113 1145 GND VDD ICV_4 $T=2904000 2784500 0 0 $X=2904000 $Y=2784500
X752 387 126 1185 1200 374 1174 1185 GND VDD ICV_4 $T=3152000 2784500 0 0 $X=3152000 $Y=2784500
X753 1224 314 388 328 377 1196 1198 GND VDD ICV_4 $T=3272000 2081500 0 0 $X=3272000 $Y=2081500
X754 1240 1293 1262 1287 1240 1246 392 GND VDD ICV_4 $T=3456000 1807500 0 0 $X=3456000 $Y=1807500
X755 152 424 152 1301 423 GND VDD ICV_5 $T=279000 618500 1 180 $X=216000 $Y=618500
X756 197 571 197 1308 573 GND VDD ICV_5 $T=759000 1341500 1 180 $X=696000 $Y=1341500
X757 202 698 i_pixel_mid[18] i_pixel_top[17] 202 GND VDD ICV_5 $T=1215000 2356500 1 180 $X=1152000 $Y=2356500
X758 754 778 759 754 803 GND VDD ICV_5 $T=1527000 2356500 1 180 $X=1464000 $Y=2356500
X759 i_pixel_top[11] 872 861 889 883 GND VDD ICV_5 $T=1895000 1474500 1 180 $X=1832000 $Y=1474500
X760 873 882 844 873 880 GND VDD ICV_5 $T=1903000 2356500 1 180 $X=1840000 $Y=2356500
X761 290 909 290 892 298 GND VDD ICV_5 $T=2007000 2501500 1 180 $X=1944000 $Y=2501500
X762 391 1258 1236 391 1279 GND VDD ICV_5 $T=3479000 1341500 1 180 $X=3416000 $Y=1341500
X763 1062 i_reset i_clock o_mode[0] GND VDD dffs_ni $T=2678000 7000 1 180 $X=2480000 $Y=7000
X764 GND i_reset i_clock 135 GND VDD dffs_ni $T=3408000 7000 0 0 $X=3408000 $Y=7000
X765 179 512 507 491 178 168 496 GND VDD ICV_6 $T=512000 2501500 0 0 $X=512000 $Y=2501500
X766 30 18 576 557 18 107 557 GND VDD ICV_6 $T=672000 7000 0 0 $X=672000 $Y=7000
X767 581 32 631 590 32 570 590 GND VDD ICV_6 $T=776000 328500 0 0 $X=776000 $Y=328500
X768 653 263 222 i_valid 232 644 648 GND VDD ICV_6 $T=1048000 328500 0 0 $X=1048000 $Y=328500
X769 84 705 733 753 705 753 706 GND VDD ICV_6 $T=1272000 2081500 0 0 $X=1272000 $Y=2081500
X770 736 237 775 748 33 726 730 GND VDD ICV_6 $T=1336000 461500 0 0 $X=1336000 $Y=461500
X771 774 254 801 782 254 762 782 GND VDD ICV_6 $T=1488000 783500 0 0 $X=1488000 $Y=783500
X772 558 825 923 272 825 272 832 GND VDD ICV_6 $T=1720000 2784500 0 0 $X=1720000 $Y=2784500
X773 881 884 905 891 62 866 891 GND VDD ICV_6 $T=1864000 1057500 0 0 $X=1864000 $Y=1057500
X774 905 908 918 912 908 897 912 GND VDD ICV_6 $T=1984000 916500 0 0 $X=1984000 $Y=916500
X775 965 968 971 i_valid 929 956 961 GND VDD ICV_6 $T=2232000 461500 0 0 $X=2232000 $Y=461500
X776 1031 973 979 969 954 973 969 GND VDD ICV_6 $T=2248000 2356500 0 0 $X=2248000 $Y=2356500
X777 362 1019 i_pixel_bot[20] 1042 1019 1042 343 GND VDD ICV_6 $T=2576000 2223500 0 0 $X=2576000 $Y=2223500
X778 360 i_pixel_bot[21] 1077 1105 1077 1105 1054 GND VDD ICV_6 $T=2792000 1807500 0 0 $X=2792000 $Y=1807500
X779 1123 367 1093 1117 1093 1117 1099 GND VDD ICV_6 $T=2848000 1057500 0 0 $X=2848000 $Y=1057500
X780 1111 362 1127 364 362 364 1057 GND VDD ICV_6 $T=2856000 2501500 0 0 $X=2856000 $Y=2501500
X781 1190 108 1139 1143 108 1143 365 GND VDD ICV_6 $T=2944000 1948500 0 0 $X=2944000 $Y=1948500
X782 1148 1133 135 1183 1133 1183 1144 GND VDD ICV_6 $T=3000000 7000 0 0 $X=3000000 $Y=7000
X783 1212 1190 1208 1210 1190 1210 380 GND VDD ICV_6 $T=3256000 1948500 0 0 $X=3256000 $Y=1948500
X784 138 i_pixel_mid[23] 1238 1256 i_pixel_mid[23] i_pixel_mid[7] 1256 GND VDD ICV_6 $T=3376000 1948500 0 0 $X=3376000 $Y=1948500
X785 162 158 433 462 GND VDD and03 $T=393500 1807500 1 180 $X=344000 $Y=1807500
X786 159 410 166 428 GND VDD and03 $T=393500 2223500 1 180 $X=344000 $Y=2223500
X787 153 552 176 562 GND VDD and03 $T=648000 461500 0 0 $X=648000 $Y=461500
X788 205 30 176 201 GND VDD and03 $T=824000 618500 0 0 $X=824000 $Y=618500
X789 729 i_pixel_bot[16] 720 758 GND VDD and03 $T=1417500 1666500 1 180 $X=1368000 $Y=1666500
X790 59 90 41 865 GND VDD and03 $T=1825500 7000 1 180 $X=1776000 $Y=7000
X791 70 91 900 1313 GND VDD and03 $T=2008000 328500 0 0 $X=2008000 $Y=328500
X792 879 i_pixel_bot[8] 288 911 GND VDD and03 $T=2056000 1948500 0 0 $X=2056000 $Y=1948500
X793 312 311 309 946 GND VDD and03 $T=2217500 1474500 1 180 $X=2168000 $Y=1474500
X794 313 331 326 96 GND VDD and03 $T=2417500 2356500 1 180 $X=2368000 $Y=2356500
X795 1138 1268 1110 1147 GND VDD and03 $T=3024000 328500 0 0 $X=3024000 $Y=328500
X796 379 1294 393 1225 GND VDD and03 $T=3376000 618500 0 0 $X=3376000 $Y=618500
X797 183 466 501 501 516 224 GND VDD ICV_7 $T=488000 1341500 0 0 $X=488000 $Y=1341500
X798 527 536 537 188 203 536 GND VDD ICV_7 $T=672000 2634500 0 0 $X=672000 $Y=2634500
X799 548 537 500 i_pixel_top[23] 558 548 GND VDD ICV_7 $T=672000 2784500 0 0 $X=672000 $Y=2784500
X800 487 517 607 665 677 487 GND VDD ICV_7 $T=904000 152500 0 0 $X=904000 $Y=152500
X801 i_pixel_mid[7] i_pixel_bot[6] 624 661 755 664 GND VDD ICV_7 $T=1024000 2634500 0 0 $X=1024000 $Y=2634500
X802 700 738 668 267 72 700 GND VDD ICV_7 $T=1184000 152500 0 0 $X=1184000 $Y=152500
X803 226 697 703 238 242 232 GND VDD ICV_7 $T=1216000 1200500 0 0 $X=1216000 $Y=1200500
X804 727 767 737 749 259 744 GND VDD ICV_7 $T=1352000 2784500 0 0 $X=1352000 $Y=2784500
X805 744 740 747 247 53 740 GND VDD ICV_7 $T=1376000 2917500 0 0 $X=1376000 $Y=2917500
X806 i_pixel_bot[10] i_pixel_top[10] 739 769 249 763 GND VDD ICV_7 $T=1432000 2223500 0 0 $X=1432000 $Y=2223500
X807 251 788 783 841 868 788 GND VDD ICV_7 $T=1536000 2634500 0 0 $X=1536000 $Y=2634500
X808 779 787 254 830 313 781 GND VDD ICV_7 $T=1568000 1341500 0 0 $X=1568000 $Y=1341500
X809 815 819 818 830 314 258 GND VDD ICV_7 $T=1664000 1200500 0 0 $X=1664000 $Y=1200500
X810 i_pixel_mid[3] i_pixel_bot[2] 804 i_pixel_mid[1] i_pixel_top[2] 873 GND VDD ICV_7 $T=1712000 2356500 0 0 $X=1712000 $Y=2356500
X811 847 851 289 255 91 862 GND VDD ICV_7 $T=1816000 328500 0 0 $X=1816000 $Y=328500
X812 836 831 927 880 869 892 GND VDD ICV_7 $T=1816000 2501500 0 0 $X=1816000 $Y=2501500
X813 871 858 62 830 309 871 GND VDD ICV_7 $T=1840000 1200500 0 0 $X=1840000 $Y=1200500
X814 852 60 274 887 87 251 GND VDD ICV_7 $T=1840000 2081500 0 0 $X=1840000 $Y=2081500
X815 i_pixel_mid[4] i_pixel_bot[3] 868 i_pixel_mid[5] i_pixel_bot[4] 859 GND VDD ICV_7 $T=1848000 2634500 0 0 $X=1848000 $Y=2634500
X816 295 273 310 943 952 908 GND VDD ICV_7 $T=2072000 1057500 0 0 $X=2072000 $Y=1057500
X817 322 331 86 i_pixel_top[3] i_pixel_top[12] 991 GND VDD ICV_7 $T=2352000 1341500 0 0 $X=2352000 $Y=1341500
X818 i_pixel_bot[5] i_pixel_top[21] 1003 i_pixel_mid[4] i_pixel_top[5] 1061 GND VDD ICV_7 $T=2376000 2501500 0 0 $X=2376000 $Y=2501500
X819 i_pixel_bot[5] i_pixel_bot[12] 1002 i_pixel_mid[19] i_pixel_bot[20] 1042 GND VDD ICV_7 $T=2448000 2223500 0 0 $X=2448000 $Y=2223500
X820 1034 1037 1024 1063 1058 350 GND VDD ICV_7 $T=2624000 1057500 0 0 $X=2624000 $Y=1057500
X821 i_pixel_bot[13] i_pixel_bot[20] 366 1109 1139 1143 GND VDD ICV_7 $T=2816000 1948500 0 0 $X=2816000 $Y=1948500
X822 i_pixel_bot[21] i_pixel_top[5] 1105 360 1151 1107 GND VDD ICV_7 $T=2848000 1666500 0 0 $X=2848000 $Y=1666500
X823 342 1126 375 1160 380 127 GND VDD ICV_7 $T=3024000 1200500 0 0 $X=3024000 $Y=1200500
X824 1154 1145 1125 1161 1185 1200 GND VDD ICV_7 $T=3024000 2784500 0 0 $X=3024000 $Y=2784500
X825 358 370 1154 i_pixel_mid[22] i_pixel_bot[23] 1174 GND VDD ICV_7 $T=3040000 2634500 0 0 $X=3040000 $Y=2634500
X826 119 1159 1214 372 1171 1262 GND VDD ICV_7 $T=3088000 1807500 0 0 $X=3088000 $Y=1807500
X827 i_pixel_bot[15] i_pixel_bot[22] 1171 1184 1208 1210 GND VDD ICV_7 $T=3128000 1948500 0 0 $X=3128000 $Y=1948500
X828 1168 1163 140 1194 383 382 GND VDD ICV_7 $T=3184000 1341500 0 0 $X=3184000 $Y=1341500
X829 637 574 600 609 564 550 534 192 609 574 GND VDD ICV_8 $T=720000 2501500 0 0 $X=720000 $Y=2501500
X830 589 215 625 624 i_pixel_bot[7] 589 203 206 624 215 GND VDD ICV_8 $T=840000 2634500 0 0 $X=840000 $Y=2634500
X831 606 629 658 651 606 617 627 651 629 635 GND VDD ICV_8 $T=944000 1474500 0 0 $X=944000 $Y=1474500
X832 594 704 670 676 832 630 634 639 676 670 GND VDD ICV_8 $T=1000000 2917500 0 0 $X=1000000 $Y=2917500
X833 80 28 706 712 i_pixel_top[18] i_pixel_top[9] 657 228 712 28 GND VDD ICV_8 $T=1072000 1948500 0 0 $X=1072000 $Y=1948500
X834 792 749 81 259 i_pixel_mid[19] i_pixel_top[18] 767 770 260 792 GND VDD ICV_8 $T=1480000 2784500 0 0 $X=1480000 $Y=2784500
X835 822 239 839 829 217 221 795 829 106 239 GND VDD ICV_8 $T=1576000 461500 0 0 $X=1576000 $Y=461500
X836 1076 345 356 1078 i_pixel_bot[7] i_pixel_bot[14] 1039 1037 1078 345 GND VDD ICV_8 $T=2568000 1666500 0 0 $X=2568000 $Y=1666500
X837 358 1043 1067 1061 1018 1025 1055 1073 1061 1043 GND VDD ICV_8 $T=2568000 2501500 0 0 $X=2568000 $Y=2501500
X838 1093 1076 351 1104 i_pixel_top[15] 1048 354 1058 1104 1076 GND VDD ICV_8 $T=2656000 1200500 0 0 $X=2656000 $Y=1200500
X839 368 1096 1116 1091 352 991 1119 1160 1091 1096 GND VDD ICV_8 $T=2760000 1341500 0 0 $X=2760000 $Y=1341500
X840 1252 139 387 390 126 1200 1205 1245 390 387 GND VDD ICV_8 $T=3272000 2784500 0 0 $X=3272000 $Y=2784500
X841 1270 1260 1249 1231 138 1219 1231 391 1231 1249 GND VDD ICV_8 $T=3352000 1666500 0 0 $X=3352000 $Y=1666500
X842 149 420 226 408 157 405 GND VDD ICV_9 $T=215000 1341500 1 180 $X=152000 $Y=1341500
X843 409 433 413 409 151 145 GND VDD ICV_9 $T=215000 1807500 1 180 $X=152000 $Y=1807500
X844 163 490 485 16 1303 1302 GND VDD ICV_9 $T=487000 618500 1 180 $X=424000 $Y=618500
X845 198 565 561 555 577 565 GND VDD ICV_9 $T=775000 1807500 1 180 $X=712000 $Y=1807500
X846 593 657 578 i_pixel_bot[15] i_pixel_top[15] 195 GND VDD ICV_9 $T=791000 1666500 1 180 $X=728000 $Y=1666500
X847 i_pixel_bot[1] i_pixel_top[17] 646 579 202 564 GND VDD ICV_9 $T=855000 2356500 1 180 $X=792000 $Y=2356500
X848 200 206 601 582 21 568 GND VDD ICV_9 $T=863000 2784500 1 180 $X=800000 $Y=2784500
X849 i_pixel_bot[9] i_pixel_top[9] 623 i_pixel_bot[2] i_pixel_bot[9] 208 GND VDD ICV_9 $T=1007000 1948500 1 180 $X=944000 $Y=1948500
X850 663 674 754 i_pixel_mid[17] i_pixel_bot[18] 674 GND VDD ICV_9 $T=1087000 2223500 1 180 $X=1024000 $Y=2223500
X851 i_pixel_bot[2] i_pixel_top[18] 731 626 739 229 GND VDD ICV_9 $T=1311000 2223500 1 180 $X=1248000 $Y=2223500
X852 764 756 60 i_pixel_bot[10] i_pixel_bot[17] 756 GND VDD ICV_9 $T=1423000 1948500 1 180 $X=1360000 $Y=1948500
X853 255 41 766 267 65 647 GND VDD ICV_9 $T=1503000 7000 1 180 $X=1440000 $Y=7000
X854 827 817 843 828 69 791 GND VDD ICV_9 $T=1671000 1807500 1 180 $X=1608000 $Y=1807500
X855 255 70 813 813 807 239 GND VDD ICV_9 $T=1703000 328500 1 180 $X=1640000 $Y=328500
X856 270 274 889 849 843 878 GND VDD ICV_9 $T=1855000 1807500 1 180 $X=1792000 $Y=1807500
X857 i_pixel_mid[18] i_pixel_mid[2] 867 893 867 852 GND VDD ICV_9 $T=1895000 2223500 1 180 $X=1832000 $Y=2223500
X858 i_pixel_mid[23] i_pixel_top[22] 272 i_pixel_mid[21] i_pixel_top[20] 259 GND VDD ICV_9 $T=2047000 2784500 1 180 $X=1984000 $Y=2784500
X859 i_pixel_bot[14] i_pixel_top[14] 301 i_pixel_bot[19] i_pixel_top[3] 69 GND VDD ICV_9 $T=2071000 1807500 1 180 $X=2008000 $Y=1807500
X860 304 315 913 913 901 300 GND VDD ICV_9 $T=2079000 1200500 1 180 $X=2016000 $Y=1200500
X861 i_pixel_top[23] i_pixel_top[14] 336 333 1059 989 GND VDD ICV_9 $T=2487000 1807500 1 180 $X=2424000 $Y=1807500
X862 i_pixel_bot[6] i_pixel_bot[13] 1049 997 1002 1016 GND VDD ICV_9 $T=2535000 2081500 1 180 $X=2472000 $Y=2081500
X863 i_pixel_top[6] i_pixel_top[15] 1163 i_pixel_bot[23] i_pixel_top[7] 1131 GND VDD ICV_9 $T=3055000 1474500 1 180 $X=2992000 $Y=1474500
X864 1232 392 1273 1218 382 1317 GND VDD ICV_9 $T=3399000 1200500 1 180 $X=3336000 $Y=1200500
X865 605 647 18 647 605 543 GND VDD ICV_10 $T=943000 7000 1 180 $X=880000 $Y=7000
X866 236 258 551 258 236 32 GND VDD ICV_10 $T=1319000 328500 1 180 $X=1256000 $Y=328500
X867 760 862 738 267 74 665 GND VDD ICV_10 $T=1375000 152500 1 180 $X=1312000 $Y=152500
X868 30 104 231 862 760 237 GND VDD ICV_10 $T=1431000 328500 1 180 $X=1368000 $Y=328500
X869 751 752 242 752 751 33 GND VDD ICV_10 $T=1455000 1200500 1 180 $X=1392000 $Y=1200500
X870 772 86 751 86 772 241 GND VDD ICV_10 $T=1471000 1341500 1 180 $X=1408000 $Y=1341500
X871 1177 371 107 371 1177 109 GND VDD ICV_10 $T=2863000 152500 1 180 $X=2800000 $Y=152500
X872 389 1182 1177 1182 389 517 GND VDD ICV_10 $T=3167000 152500 1 180 $X=3104000 $Y=152500
X873 134 1213 389 1213 134 101 GND VDD ICV_10 $T=3343000 461500 1 180 $X=3280000 $Y=461500
X874 436 162 466 9 164 GND VDD and04 $T=360000 1666500 0 0 $X=360000 $Y=1666500
X875 151 147 157 428 463 GND VDD and04 $T=400000 1807500 0 0 $X=400000 $Y=1807500
X876 743 59 39 61 761 GND VDD and04 $T=1481500 152500 1 180 $X=1424000 $Y=152500
X877 72 65 74 1313 907 GND VDD and04 $T=2016000 152500 0 0 $X=2016000 $Y=152500
X878 955 312 315 269 858 GND VDD and04 $T=2104000 1341500 0 0 $X=2104000 $Y=1341500
X879 334 314 376 96 330 GND VDD and04 $T=2360000 1807500 0 0 $X=2360000 $Y=1807500
X880 369 1138 118 98 1164 GND VDD and04 $T=3065500 618500 1 180 $X=3008000 $Y=618500
X881 1209 128 381 1225 1195 GND VDD and04 $T=3248000 618500 0 0 $X=3248000 $Y=618500
X882 411 419 152 412 153 VDD GND aoi22 $T=257000 328500 1 180 $X=208000 $Y=328500
X883 456 169 16 479 153 VDD GND aoi22 $T=433000 461500 1 180 $X=384000 $Y=461500
X884 480 477 152 543 472 VDD GND aoi22 $T=513000 152500 1 180 $X=464000 $Y=152500
X885 186 169 163 518 196 VDD GND aoi22 $T=641000 618500 1 180 $X=592000 $Y=618500
X886 560 169 189 553 196 VDD GND aoi22 $T=793000 783500 1 180 $X=744000 $Y=783500
X887 575 29 197 556 196 VDD GND aoi22 $T=809000 1057500 1 180 $X=760000 $Y=1057500
X888 587 194 199 31 575 VDD GND aoi22 $T=792000 916500 0 0 $X=792000 $Y=916500
X889 194 29 209 603 196 VDD GND aoi22 $T=865000 1057500 1 180 $X=816000 $Y=1057500
X890 595 234 189 217 612 VDD GND aoi22 $T=913000 783500 1 180 $X=864000 $Y=783500
X891 604 20 226 42 196 VDD GND aoi22 $T=953000 1057500 1 180 $X=904000 $Y=1057500
X892 1309 234 16 668 612 VDD GND aoi22 $T=1009000 618500 1 180 $X=960000 $Y=618500
X893 622 20 210 216 196 VDD GND aoi22 $T=1009000 1057500 1 180 $X=960000 $Y=1057500
X894 682 234 210 239 612 VDD GND aoi22 $T=1177000 783500 1 180 $X=1128000 $Y=783500
X895 734 234 209 833 612 VDD GND aoi22 $T=1409000 1057500 1 180 $X=1360000 $Y=1057500
X896 769 739 626 733 i_pixel_top[10] VDD GND aoi22 $T=1425000 2223500 1 180 $X=1376000 $Y=2223500
X897 836 731 724 243 i_pixel_bot[2] VDD GND aoi22 $T=1376000 2356500 0 0 $X=1376000 $Y=2356500
X898 828 40 768 784 i_pixel_top[2] VDD GND aoi22 $T=1569000 1807500 1 180 $X=1520000 $Y=1807500
X899 967 867 893 899 i_pixel_mid[2] VDD GND aoi22 $T=2009000 2223500 1 180 $X=1960000 $Y=2223500
X900 76 301 906 103 i_pixel_top[14] VDD GND aoi22 $T=2081000 2081500 1 180 $X=2032000 $Y=2081500
X901 932 87 887 94 i_pixel_top[12] VDD GND aoi22 $T=2313000 2081500 1 180 $X=2264000 $Y=2081500
X902 1047 966 982 923 i_pixel_bot[6] VDD GND aoi22 $T=2296000 2784500 0 0 $X=2296000 $Y=2784500
X903 994 985 987 81 i_pixel_bot[4] VDD GND aoi22 $T=2376000 2634500 0 0 $X=2376000 $Y=2634500
X904 1077 1059 333 1112 i_pixel_top[4] VDD GND aoi22 $T=2785000 1807500 1 180 $X=2736000 $Y=1807500
X905 1152 1075 1079 1082 i_pixel_mid[4] VDD GND aoi22 $T=2784000 2081500 0 0 $X=2784000 $Y=2081500
X906 1122 1151 360 1157 i_pixel_top[6] VDD GND aoi22 $T=3025000 1666500 1 180 $X=2976000 $Y=1666500
X907 1238 1196 377 1187 i_pixel_mid[6] VDD GND aoi22 $T=3216000 2081500 0 0 $X=3216000 $Y=2081500
X908 507 188 527 536 188 567 491 507 491 171 GND VDD ICV_11 $T=551000 2634500 1 180 $X=488000 $Y=2634500
X909 213 561 596 617 578 561 617 213 679 193 GND VDD ICV_11 $T=791000 1474500 1 180 $X=728000 $Y=1474500
X910 75 227 786 250 i_pixel_top[19] i_pixel_top[10] 250 227 250 742 GND VDD ICV_11 $T=1471000 1474500 1 180 $X=1408000 $Y=1474500
X911 100 919 939 914 919 914 954 i_pixel_mid[2] i_pixel_top[3] 914 GND VDD ICV_11 $T=2063000 2356500 1 180 $X=2000000 $Y=2356500
X912 1019 79 949 925 79 925 308 i_pixel_mid[18] i_pixel_bot[19] 925 GND VDD ICV_11 $T=2111000 2223500 1 180 $X=2048000 $Y=2223500
X913 99 80 957 980 84 316 957 i_pixel_bot[4] i_pixel_bot[11] 316 GND VDD ICV_11 $T=2175000 1948500 1 180 $X=2112000 $Y=1948500
X914 1009 305 993 976 305 976 983 i_pixel_top[21] i_pixel_top[12] 976 GND VDD ICV_11 $T=2311000 1200500 1 180 $X=2248000 $Y=1200500
X915 1043 100 i_pixel_top[4] 1004 100 1004 1018 i_pixel_mid[3] i_pixel_top[4] 1004 GND VDD ICV_11 $T=2487000 2356500 1 180 $X=2424000 $Y=2356500
X916 385 1178 1192 1173 1178 1173 1193 i_pixel_mid[6] i_pixel_top[7] 1173 GND VDD ICV_11 $T=3159000 2501500 1 180 $X=3096000 $Y=2501500
X917 1293 1212 1214 1199 1212 1199 383 1198 1214 1199 GND VDD ICV_11 $T=3279000 1807500 1 180 $X=3216000 $Y=1807500
X918 465 147 469 125 409 159 161 GND VDD ICV_12 $T=407000 1948500 1 180 $X=344000 $Y=1948500
X919 481 514 478 471 514 471 461 GND VDD ICV_12 $T=455000 1057500 1 180 $X=392000 $Y=1057500
X920 178 513 503 500 503 500 173 GND VDD ICV_12 $T=583000 2784500 1 180 $X=520000 $Y=2784500
X921 592 487 684 607 543 109 566 GND VDD ICV_12 $T=847000 152500 1 180 $X=784000 $Y=152500
X922 661 667 637 690 637 690 550 GND VDD ICV_12 $T=1079000 2501500 1 180 $X=1016000 $Y=2501500
X923 893 i_pixel_mid[17] 816 797 i_pixel_mid[17] i_pixel_mid[1] 797 GND VDD ICV_12 $T=1623000 2223500 1 180 $X=1560000 $Y=2223500
X924 987 i_pixel_top[19] 836 831 i_pixel_bot[3] i_pixel_top[19] 831 GND VDD ICV_12 $T=1759000 2501500 1 180 $X=1696000 $Y=2501500
X925 305 75 i_pixel_top[11] 926 i_pixel_top[20] i_pixel_top[11] 926 GND VDD ICV_12 $T=2047000 1474500 1 180 $X=1984000 $Y=1474500
X926 1013 941 308 953 927 308 953 GND VDD ICV_12 $T=2159000 2501500 1 180 $X=2096000 $Y=2501500
X927 329 970 981 964 958 970 964 GND VDD ICV_12 $T=2287000 1474500 1 180 $X=2224000 $Y=1474500
X928 1079 i_pixel_mid[19] 967 984 967 984 977 GND VDD ICV_12 $T=2327000 2223500 1 180 $X=2264000 $Y=2223500
X929 108 92 88 998 977 88 998 GND VDD ICV_12 $T=2359000 1948500 1 180 $X=2296000 $Y=1948500
X930 1026 338 329 975 983 338 975 GND VDD ICV_12 $T=2383000 1057500 1 180 $X=2320000 $Y=1057500
X931 1012 1008 337 i_valid 999 1102 992 GND VDD ICV_12 $T=2503000 618500 1 180 $X=2440000 $Y=618500
X932 339 1009 i_pixel_top[13] 1022 i_pixel_top[22] i_pixel_top[13] 1022 GND VDD ICV_12 $T=2503000 1057500 1 180 $X=2440000 $Y=1057500
X933 342 335 1315 1023 1001 335 1023 GND VDD ICV_12 $T=2511000 1666500 1 180 $X=2448000 $Y=1666500
X934 353 1037 1026 1024 1026 1024 337 GND VDD ICV_12 $T=2583000 916500 1 180 $X=2520000 $Y=916500
X935 1149 63 i_pixel_bot[19] 1066 i_pixel_bot[12] i_pixel_bot[19] 1066 GND VDD ICV_12 $T=2663000 1948500 1 180 $X=2600000 $Y=1948500
X936 1086 1058 353 350 1046 1103 349 GND VDD ICV_12 $T=2703000 916500 1 180 $X=2640000 $Y=916500
X937 1129 1087 1088 359 1073 1087 359 GND VDD ICV_12 $T=2799000 2634500 1 180 $X=2736000 $Y=2634500
X938 372 119 i_pixel_bot[21] 1159 i_pixel_bot[14] i_pixel_bot[21] 1159 GND VDD ICV_12 $T=3031000 1807500 1 180 $X=2968000 $Y=1807500
X939 1178 358 i_pixel_top[6] 370 i_pixel_mid[5] i_pixel_top[6] 370 GND VDD ICV_12 $T=3039000 2501500 1 180 $X=2976000 $Y=2501500
X940 377 i_pixel_mid[21] 1152 1150 i_pixel_mid[21] i_pixel_mid[5] 1150 GND VDD ICV_12 $T=3063000 2081500 1 180 $X=3000000 $Y=2081500
X941 404 o_edge 167 411 1300 GND VDD nand04 $T=152000 328500 0 0 $X=152000 $Y=328500
X942 463 493 462 466 9 GND VDD nand04 $T=424000 1666500 0 0 $X=424000 $Y=1666500
X943 907 864 865 39 61 GND VDD nand04 $T=1872000 7000 0 0 $X=1872000 $Y=7000
X944 330 1314 946 315 269 GND VDD nand04 $T=2200000 1341500 0 0 $X=2200000 $Y=1341500
X945 1056 104 1027 1044 1060 GND VDD nand04 $T=2641000 461500 1 180 $X=2592000 $Y=461500
X946 1195 1134 1147 118 98 GND VDD nand04 $T=3000000 461500 0 0 $X=3000000 $Y=461500
X947 711 715 225 721 737 664 21 219 721 225 GND VDD ICV_13 $T=1104000 2784500 0 0 $X=1104000 $Y=2784500
X948 841 253 811 804 763 780 755 780 804 253 GND VDD ICV_13 $T=1512000 2501500 0 0 $X=1512000 $Y=2501500
X949 290 790 1311 264 i_pixel_bot[11] i_pixel_bot[18] 257 264 790 842 GND VDD ICV_13 $T=1608000 2081500 0 0 $X=1608000 $Y=2081500
X950 898 878 902 273 830 311 815 273 878 857 GND VDD ICV_13 $T=1760000 1341500 0 0 $X=1760000 $Y=1341500
X951 1053 1013 343 1017 987 985 1011 1017 343 1011 GND VDD ICV_13 $T=2432000 2634500 0 0 $X=2432000 $Y=2634500
X952 139 i_pixel_top[23] 1047 1041 i_pixel_bot[7] i_pixel_top[23] 1041 1035 1057 1036 GND VDD ICV_13 $T=2536000 2784500 0 0 $X=2536000 $Y=2784500
X953 126 1101 1097 1113 1047 1041 1161 1113 1097 114 GND VDD ICV_13 $T=2720000 2784500 0 0 $X=2720000 $Y=2784500
X954 367 i_pixel_bot[23] 1122 1131 i_pixel_top[5] i_pixel_top[14] 1128 1100 1131 1122 GND VDD ICV_13 $T=2808000 1474500 0 0 $X=2808000 $Y=1474500
X955 1135 1141 1123 1120 1086 1070 361 1103 1120 1123 GND VDD ICV_13 $T=2816000 916500 0 0 $X=2816000 $Y=916500
X956 1142 365 342 1126 1100 351 1104 1126 365 1119 GND VDD ICV_13 $T=2840000 1200500 0 0 $X=2840000 $Y=1200500
X957 8 1307 495 540 GND VDD mux21_ni $T=664000 1474500 0 0 $X=664000 $Y=1474500
X958 572 581 14 591 GND VDD mux21_ni $T=808000 461500 0 0 $X=808000 $Y=461500
X959 123 800 261 856 GND VDD mux21_ni $T=1670000 783500 1 180 $X=1608000 $Y=783500
X960 809 61 98 931 GND VDD mux21_ni $T=2206000 783500 1 180 $X=2144000 $Y=783500
X961 123 951 319 986 GND VDD mux21_ni $T=2270000 783500 1 180 $X=2208000 $Y=783500
X962 129 268 320 978 GND VDD mux21_ni $T=2326000 916500 1 180 $X=2264000 $Y=916500
X963 344 1165 o_mode[0] 1062 GND VDD mux21_ni $T=2680000 7000 0 0 $X=2680000 $Y=7000
X964 355 i_valid 1114 1089 GND VDD mux21_ni $T=2806000 7000 1 180 $X=2744000 $Y=7000
X965 VDD 67 324 280 GND VDD latchr $T=1981000 783500 1 180 $X=1896000 $Y=783500
X966 VDD 306 324 936 GND VDD latchr $T=2112000 152500 0 0 $X=2112000 $Y=152500
X967 VDD 960 324 1289 GND VDD latchr $T=2248000 618500 0 0 $X=2248000 $Y=618500
X968 544 528 1307 9 i_valid GND VDD oai22 $T=672000 1666500 0 0 $X=672000 $Y=1666500
X969 240 244 800 61 i_valid GND VDD oai22 $T=1481000 783500 1 180 $X=1432000 $Y=783500
X970 834 837 268 269 i_valid GND VDD oai22 $T=1776000 1474500 0 0 $X=1776000 $Y=1474500
X971 307 318 951 98 i_valid GND VDD oai22 $T=2208000 916500 0 0 $X=2208000 $Y=916500
X972 474 461 167 509 GND VDD oai21 $T=465000 916500 1 180 $X=424000 $Y=916500
X973 i_pixel_mid[16] 547 526 191 GND VDD oai21 $T=705000 2081500 1 180 $X=664000 $Y=2081500
X974 579 i_pixel_mid[17] 542 i_pixel_top[16] GND VDD oai21 $T=745000 2356500 1 180 $X=704000 $Y=2356500
X975 593 i_pixel_top[17] 635 i_pixel_top[8] GND VDD oai21 $T=896000 1666500 0 0 $X=896000 $Y=1666500
X976 598 i_pixel_bot[1] 207 i_pixel_bot[8] GND VDD oai21 $T=937000 1948500 1 180 $X=896000 $Y=1948500
X977 20 52 640 224 GND VDD oai21 $T=1057000 916500 1 180 $X=1016000 $Y=916500
X978 640 218 669 672 GND VDD oai21 $T=1064000 916500 0 0 $X=1064000 $Y=916500
X979 663 i_pixel_mid[16] 654 i_pixel_bot[17] GND VDD oai21 $T=1145000 2081500 1 180 $X=1104000 $Y=2081500
X980 713 218 693 672 GND VDD oai21 $T=1128000 1057500 0 0 $X=1128000 $Y=1057500
X981 692 i_pixel_mid[1] 600 i_pixel_bot[0] GND VDD oai21 $T=1193000 2634500 1 180 $X=1152000 $Y=2634500
X982 686 741 27 683 GND VDD oai21 $T=1217000 916500 1 180 $X=1176000 $Y=916500
X983 713 734 707 718 GND VDD oai21 $T=1321000 1057500 1 180 $X=1280000 $Y=1057500
X984 i_pixel_top[16] 719 666 235 GND VDD oai21 $T=1353000 1474500 1 180 $X=1312000 $Y=1474500
X985 i_pixel_top[0] 750 826 758 GND VDD oai21 $T=1472000 1666500 0 0 $X=1472000 $Y=1666500
X986 764 i_pixel_bot[9] 817 i_pixel_bot[16] GND VDD oai21 $T=1520000 1948500 0 0 $X=1520000 $Y=1948500
X987 824 i_pixel_top[0] 857 i_pixel_top[9] GND VDD oai21 $T=1664000 1474500 0 0 $X=1664000 $Y=1474500
X988 12 776 921 821 GND VDD oai21 $T=1672000 618500 0 0 $X=1672000 $Y=618500
X989 844 i_pixel_mid[0] 842 i_pixel_top[1] GND VDD oai21 $T=1792000 2081500 0 0 $X=1792000 $Y=2081500
X990 i_pixel_top[8] 916 295 911 GND VDD oai21 $T=2057000 1666500 1 180 $X=2016000 $Y=1666500
X991 320 283 935 931 GND VDD oai21 $T=2160000 916500 0 0 $X=2160000 $Y=916500
X992 107 177 18 VDD GND nor02 $T=552000 152500 0 0 $X=552000 $Y=152500
X993 177 559 231 VDD GND nor02 $T=704000 461500 0 0 $X=704000 $Y=461500
X994 549 570 231 VDD GND nor02 $T=736000 328500 0 0 $X=736000 $Y=328500
X995 608 644 231 VDD GND nor02 $T=952000 328500 0 0 $X=952000 $Y=328500
X996 660 762 231 VDD GND nor02 $T=1128000 618500 0 0 $X=1128000 $Y=618500
X997 656 726 231 VDD GND nor02 $T=1240000 461500 0 0 $X=1240000 $Y=461500
X998 714 735 231 VDD GND nor02 $T=1312000 618500 0 0 $X=1312000 $Y=618500
X999 49 793 283 VDD GND nor02 $T=1600000 916500 0 0 $X=1600000 $Y=916500
X1000 54 805 283 VDD GND nor02 $T=1673000 1057500 1 180 $X=1640000 $Y=1057500
X1001 283 866 840 VDD GND nor02 $T=1825000 1057500 1 180 $X=1792000 $Y=1057500
X1002 886 897 283 VDD GND nor02 $T=1944000 916500 0 0 $X=1944000 $Y=916500
X1003 903 920 283 VDD GND nor02 $T=2040000 783500 0 0 $X=2040000 $Y=783500
X1004 344 o_mode[1] 438 VDD GND or02 $T=344000 1057500 0 0 $X=344000 $Y=1057500
X1005 i_pixel_top[8] 602 597 VDD GND or02 $T=888000 2223500 0 0 $X=888000 $Y=2223500
X1006 688 i_pixel_top[0] 655 VDD GND or02 $T=1161000 1666500 1 180 $X=1120000 $Y=1666500
X1007 746 i_pixel_bot[0] 720 VDD GND or02 $T=1377000 1807500 1 180 $X=1336000 $Y=1807500
X1008 281 i_pixel_mid[0] 288 VDD GND or02 $T=1960000 1948500 0 0 $X=1960000 $Y=1948500
X1009 619 i_pixel_bot[8] i_pixel_bot[1] 705 i_pixel_bot[9] i_pixel_bot[2] VDD GND aoi32 $T=993000 2081500 1 180 $X=936000 $Y=2081500
X1010 20 52 659 686 669 707 VDD GND aoi32 $T=1112000 916500 0 0 $X=1112000 $Y=916500
X1011 675 i_pixel_top[8] i_pixel_top[17] 227 i_pixel_top[9] i_pixel_top[18] VDD GND aoi32 $T=1160000 1807500 0 0 $X=1160000 $Y=1807500
X1012 695 i_pixel_bot[17] i_pixel_mid[16] 79 i_pixel_bot[18] i_pixel_mid[17] VDD GND aoi32 $T=1241000 2223500 1 180 $X=1184000 $Y=2223500
X1013 698 i_pixel_top[16] i_pixel_mid[17] 727 i_pixel_top[17] i_pixel_mid[18] VDD GND aoi32 $T=1248000 2356500 0 0 $X=1248000 $Y=2356500
X1014 732 i_pixel_bot[0] i_pixel_mid[1] 253 i_pixel_bot[1] i_pixel_mid[2] VDD GND aoi32 $T=1392000 2501500 0 0 $X=1392000 $Y=2501500
X1015 777 i_pixel_bot[16] i_pixel_bot[9] 820 i_pixel_bot[17] i_pixel_bot[10] VDD GND aoi32 $T=1568000 1948500 0 0 $X=1568000 $Y=1948500
X1016 808 i_pixel_top[9] i_pixel_top[0] 64 i_pixel_top[10] i_pixel_top[1] VDD GND aoi32 $T=1664000 1666500 0 0 $X=1664000 $Y=1666500
X1017 882 i_pixel_top[1] i_pixel_mid[0] 919 i_pixel_top[2] i_pixel_mid[1] VDD GND aoi32 $T=1936000 2356500 0 0 $X=1936000 $Y=2356500
X1018 585 554 i_pixel_mid[0] 597 VDD GND nand03 $T=752000 2223500 0 0 $X=752000 $Y=2223500
X1019 585 574 i_pixel_mid[0] 597 VDD GND nand03 $T=800000 2223500 0 0 $X=800000 $Y=2223500
X1020 691 211 i_pixel_bot[0] 655 VDD GND nand03 $T=1113000 1666500 1 180 $X=1072000 $Y=1666500
X1021 691 717 i_pixel_bot[0] 655 VDD GND nand03 $T=1281000 1666500 1 180 $X=1240000 $Y=1666500
X1022 729 701 i_pixel_bot[16] 720 VDD GND nand03 $T=1329000 1807500 1 180 $X=1288000 $Y=1807500
X1023 879 849 i_pixel_bot[8] 288 VDD GND nand03 $T=1913000 1948500 1 180 $X=1872000 $Y=1948500
X1024 447 551 505 437 419 107 GND VDD aoi221 $T=360000 328500 0 0 $X=360000 $Y=328500
X1025 508 232 505 185 169 517 GND VDD aoi221 $T=641000 328500 1 180 $X=576000 $Y=328500
X1026 515 32 505 165 169 109 GND VDD aoi221 $T=657000 152500 1 180 $X=592000 $Y=152500
X1027 621 33 220 498 169 101 GND VDD aoi221 $T=985000 783500 1 180 $X=920000 $Y=783500
X1028 638 254 220 199 29 221 GND VDD aoi221 $T=1056000 783500 0 0 $X=1056000 $Y=783500
X1029 693 34 699 683 29 224 GND VDD aoi221 $T=1241000 1057500 1 180 $X=1176000 $Y=1057500
X1030 694 248 220 31 29 106 GND VDD aoi221 $T=1224000 916500 0 0 $X=1224000 $Y=916500
X1031 709 241 220 546 20 136 GND VDD aoi221 $T=1296000 916500 0 0 $X=1296000 $Y=916500
X1032 153 620 154 419 422 GND VDD ao22 $T=264000 328500 0 0 $X=264000 $Y=328500
X1033 472 18 146 477 447 GND VDD ao22 $T=457500 152500 1 180 $X=400000 $Y=152500
X1034 472 487 154 477 508 GND VDD ao22 $T=521500 328500 1 180 $X=464000 $Y=328500
X1035 612 237 163 234 709 GND VDD ao22 $T=1216000 783500 0 0 $X=1216000 $Y=783500
X1036 477 201 GND VDD buf02 $T=513500 461500 1 180 $X=480000 $Y=461500
X1037 505 562 GND VDD buf02 $T=608000 461500 0 0 $X=608000 $Y=461500
X1038 234 201 GND VDD buf02 $T=817500 618500 1 180 $X=784000 $Y=618500
X1039 220 562 GND VDD buf02 $T=937500 461500 1 180 $X=904000 $Y=461500
.ENDS
***************************************
